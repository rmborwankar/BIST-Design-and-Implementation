
//Verilog file of module fourFunc


`timescale 1 ns / 1ns

module fourFunc_net(clk,
rst,
start,
func,
x,
busy,
resultIPart,
resultFPart);
	input	clk;
	input	rst;
	input	start;
input [0:1]func;
input [0:7]x;
	output 	busy;
output [0:1]resultIPart;
output [0:7]resultFPart;
wire
fourFunc_wire_1,
fourFunc_wire_2,
fourFunc_wire_3,
fourFunc_wire_4,
fourFunc_wire_5,
fourFunc_wire_6,
fourFunc_wire_7,
fourFunc_wire_8,
fourFunc_wire_9,
fourFunc_wire_10,
fourFunc_wire_11,
fourFunc_wire_12,
fourFunc_wire_13,
fourFunc_wire_14,
fourFunc_wire_15,
fourFunc_wire_16,
fourFunc_wire_17,
fourFunc_wire_18,
fourFunc_wire_19,
fourFunc_wire_20,
fourFunc_wire_21,
fourFunc_wire_22,
fourFunc_wire_23,
fourFunc_wire_24,
fourFunc_wire_25,
fourFunc_wire_26,
fourFunc_wire_27,
fourFunc_wire_28,
fourFunc_wire_29,
fourFunc_wire_30,
fourFunc_wire_31,
fourFunc_wire_32,
fourFunc_wire_33,
fourFunc_wire_34,
fourFunc_wire_35,
fourFunc_wire_36,
fourFunc_wire_37,
fourFunc_wire_38,
fourFunc_wire_39,
fourFunc_wire_40,
fourFunc_wire_41,
fourFunc_wire_42,
fourFunc_wire_43,
fourFunc_wire_44,
fourFunc_wire_45,
fourFunc_wire_46,
fourFunc_wire_47,
fourFunc_wire_48,
fourFunc_wire_49,
fourFunc_wire_50,
fourFunc_wire_51,
fourFunc_wire_52,
fourFunc_wire_53,
fourFunc_wire_54,
fourFunc_wire_55,
fourFunc_wire_56,
fourFunc_wire_57,
fourFunc_wire_58,
fourFunc_wire_59,
fourFunc_wire_60,
fourFunc_wire_61,
fourFunc_wire_62,
fourFunc_wire_63,
fourFunc_wire_64,
fourFunc_wire_65,
fourFunc_wire_66,
fourFunc_wire_67,
fourFunc_wire_68,
fourFunc_wire_69,
fourFunc_wire_70,
fourFunc_wire_71,
fourFunc_wire_72,
fourFunc_wire_73,
fourFunc_wire_74,
fourFunc_wire_75,
fourFunc_wire_76,
fourFunc_wire_77,
fourFunc_wire_78,
fourFunc_wire_79,
fourFunc_wire_80,
fourFunc_wire_81,
fourFunc_wire_82,
fourFunc_wire_83,
fourFunc_wire_84,
fourFunc_wire_85,
fourFunc_wire_86,
fourFunc_wire_87,
fourFunc_wire_88,
fourFunc_wire_89,
fourFunc_wire_90,
fourFunc_wire_91,
fourFunc_wire_92,
fourFunc_wire_93,
fourFunc_wire_94,
fourFunc_wire_95,
fourFunc_wire_96,
fourFunc_wire_97,
fourFunc_wire_98,
fourFunc_wire_99,
fourFunc_wire_100,
fourFunc_wire_101,
fourFunc_wire_102,
fourFunc_wire_103,
fourFunc_wire_104,
fourFunc_wire_105,
fourFunc_wire_106,
fourFunc_wire_107,
fourFunc_wire_108,
fourFunc_wire_109,
fourFunc_wire_110,
fourFunc_wire_111,
fourFunc_wire_112,
fourFunc_wire_113,
fourFunc_wire_114,
fourFunc_wire_115,
fourFunc_wire_116,
fourFunc_wire_117,
fourFunc_wire_118,
fourFunc_wire_119,
fourFunc_wire_120,
fourFunc_wire_121,
fourFunc_wire_122,
fourFunc_wire_123,
fourFunc_wire_124,
fourFunc_wire_125,
fourFunc_wire_126,
fourFunc_wire_127,
fourFunc_wire_128,
fourFunc_wire_129,
fourFunc_wire_130,
fourFunc_wire_131,
fourFunc_wire_132,
fourFunc_wire_133,
fourFunc_wire_134,
fourFunc_wire_135,
fourFunc_wire_136,
fourFunc_wire_137,
fourFunc_wire_138,
fourFunc_wire_139,
fourFunc_wire_140,
fourFunc_wire_141,
fourFunc_wire_142,
fourFunc_wire_143,
fourFunc_wire_144,
fourFunc_wire_145,
fourFunc_wire_146,
fourFunc_wire_147,
fourFunc_wire_148,
fourFunc_wire_149,
fourFunc_wire_150,
fourFunc_wire_151,
fourFunc_wire_152,
fourFunc_wire_153,
fourFunc_wire_154,
fourFunc_wire_155,
fourFunc_wire_156,
fourFunc_wire_157,
fourFunc_wire_158,
fourFunc_wire_159,
fourFunc_wire_160,
fourFunc_wire_161,
fourFunc_wire_162,
fourFunc_wire_163,
fourFunc_wire_164,
fourFunc_wire_165,
fourFunc_wire_166,
fourFunc_wire_167,
fourFunc_wire_168,
fourFunc_wire_169,
fourFunc_wire_170,
fourFunc_wire_171,
fourFunc_wire_172,
fourFunc_wire_173,
fourFunc_wire_174,
fourFunc_wire_175,
fourFunc_wire_176,
fourFunc_wire_177,
fourFunc_wire_178,
fourFunc_wire_179,
fourFunc_wire_180,
fourFunc_wire_181,
fourFunc_wire_182,
fourFunc_wire_183,
fourFunc_wire_184,
fourFunc_wire_185,
fourFunc_wire_186,
fourFunc_wire_187,
fourFunc_wire_188,
fourFunc_wire_189,
fourFunc_wire_190,
fourFunc_wire_191,
fourFunc_wire_192,
fourFunc_wire_193,
fourFunc_wire_194,
fourFunc_wire_195,
fourFunc_wire_196,
fourFunc_wire_197,
fourFunc_wire_198,
fourFunc_wire_199,
fourFunc_wire_200,
fourFunc_wire_201,
fourFunc_wire_202,
fourFunc_wire_203,
fourFunc_wire_204,
fourFunc_wire_205,
fourFunc_wire_206,
fourFunc_wire_207,
fourFunc_wire_208,
fourFunc_wire_209,
fourFunc_wire_210,
fourFunc_wire_211,
fourFunc_wire_212,
fourFunc_wire_213,
fourFunc_wire_214,
fourFunc_wire_215,
fourFunc_wire_216,
fourFunc_wire_217,
fourFunc_wire_218,
fourFunc_wire_219,
fourFunc_wire_220,
fourFunc_wire_221,
fourFunc_wire_222,
fourFunc_wire_223,
fourFunc_wire_224,
fourFunc_wire_225,
fourFunc_wire_226,
fourFunc_wire_227,
fourFunc_wire_228,
fourFunc_wire_229,
fourFunc_wire_230,
fourFunc_wire_231,
fourFunc_wire_232,
fourFunc_wire_233,
fourFunc_wire_234,
fourFunc_wire_235,
fourFunc_wire_236,
fourFunc_wire_237,
fourFunc_wire_238,
fourFunc_wire_239,
fourFunc_wire_240,
fourFunc_wire_241,
fourFunc_wire_242,
fourFunc_wire_243,
fourFunc_wire_244,
fourFunc_wire_245,
fourFunc_wire_246,
fourFunc_wire_247,
fourFunc_wire_248,
fourFunc_wire_249,
fourFunc_wire_250,
fourFunc_wire_251,
fourFunc_wire_252,
fourFunc_wire_253,
fourFunc_wire_254,
fourFunc_wire_255,
fourFunc_wire_256,
fourFunc_wire_257,
fourFunc_wire_258,
fourFunc_wire_259,
fourFunc_wire_260,
fourFunc_wire_261,
fourFunc_wire_262,
fourFunc_wire_263,
fourFunc_wire_264,
fourFunc_wire_265,
fourFunc_wire_266,
fourFunc_wire_267,
fourFunc_wire_268,
fourFunc_wire_269,
fourFunc_wire_270,
fourFunc_wire_271,
fourFunc_wire_272,
fourFunc_wire_273,
fourFunc_wire_274,
fourFunc_wire_275,
fourFunc_wire_276,
fourFunc_wire_277,
fourFunc_wire_278,
fourFunc_wire_279,
fourFunc_wire_280,
fourFunc_wire_281,
fourFunc_wire_282,
fourFunc_wire_283,
fourFunc_wire_284,
fourFunc_wire_285,
fourFunc_wire_286,
fourFunc_wire_287,
fourFunc_wire_288,
fourFunc_wire_289,
fourFunc_wire_290,
fourFunc_wire_291,
fourFunc_wire_292,
fourFunc_wire_293,
fourFunc_wire_294,
fourFunc_wire_295,
fourFunc_wire_296,
fourFunc_wire_297,
fourFunc_wire_298,
fourFunc_wire_299,
fourFunc_wire_300,
fourFunc_wire_301,
fourFunc_wire_302,
fourFunc_wire_303,
fourFunc_wire_304,
fourFunc_wire_305,
fourFunc_wire_306,
fourFunc_wire_307,
fourFunc_wire_308,
fourFunc_wire_309,
fourFunc_wire_310,
fourFunc_wire_311,
fourFunc_wire_312,
fourFunc_wire_313,
fourFunc_wire_314,
fourFunc_wire_315,
fourFunc_wire_316,
fourFunc_wire_317,
fourFunc_wire_318,
fourFunc_wire_319,
fourFunc_wire_320,
fourFunc_wire_321,
fourFunc_wire_322,
fourFunc_wire_323,
fourFunc_wire_324,
fourFunc_wire_325,
fourFunc_wire_326,
fourFunc_wire_327,
fourFunc_wire_328,
fourFunc_wire_329,
fourFunc_wire_330,
fourFunc_wire_331,
fourFunc_wire_332,
fourFunc_wire_333,
fourFunc_wire_334,
fourFunc_wire_335,
fourFunc_wire_336,
fourFunc_wire_337,
fourFunc_wire_338,
fourFunc_wire_339,
fourFunc_wire_340,
fourFunc_wire_341,
fourFunc_wire_342,
fourFunc_wire_343,
fourFunc_wire_344,
fourFunc_wire_345,
fourFunc_wire_346,
fourFunc_wire_347,
fourFunc_wire_348,
fourFunc_wire_349,
fourFunc_wire_350,
fourFunc_wire_351,
fourFunc_wire_352,
fourFunc_wire_353,
fourFunc_wire_354,
fourFunc_wire_355,
fourFunc_wire_356,
fourFunc_wire_357,
fourFunc_wire_358,
fourFunc_wire_359,
fourFunc_wire_360,
fourFunc_wire_361,
fourFunc_wire_362,
fourFunc_wire_363,
fourFunc_wire_364,
fourFunc_wire_365,
fourFunc_wire_366,
fourFunc_wire_367,
fourFunc_wire_368,
fourFunc_wire_369,
fourFunc_wire_370,
fourFunc_wire_371,
fourFunc_wire_372,
fourFunc_wire_373,
fourFunc_wire_374,
fourFunc_wire_375,
fourFunc_wire_376,
fourFunc_wire_377,
fourFunc_wire_378,
fourFunc_wire_379,
fourFunc_wire_380,
fourFunc_wire_381,
fourFunc_wire_382,
fourFunc_wire_383,
fourFunc_wire_384,
fourFunc_wire_385,
fourFunc_wire_386,
fourFunc_wire_387,
fourFunc_wire_388,
fourFunc_wire_389,
fourFunc_wire_390,
fourFunc_wire_391,
fourFunc_wire_392,
fourFunc_wire_393,
fourFunc_wire_394,
fourFunc_wire_395,
fourFunc_wire_396,
fourFunc_wire_397,
fourFunc_wire_398,
fourFunc_wire_399,
fourFunc_wire_400,
fourFunc_wire_401,
fourFunc_wire_402,
fourFunc_wire_403,
fourFunc_wire_404,
fourFunc_wire_405,
fourFunc_wire_406,
fourFunc_wire_407,
fourFunc_wire_408,
fourFunc_wire_409,
fourFunc_wire_410,
fourFunc_wire_411,
fourFunc_wire_412,
fourFunc_wire_413,
fourFunc_wire_414,
fourFunc_wire_415,
fourFunc_wire_416,
fourFunc_wire_417,
fourFunc_wire_418,
fourFunc_wire_419,
fourFunc_wire_420,
fourFunc_wire_421,
fourFunc_wire_422,
fourFunc_wire_423,
fourFunc_wire_424,
fourFunc_wire_425,
fourFunc_wire_426,
fourFunc_wire_427,
fourFunc_wire_428,
fourFunc_wire_429,
fourFunc_wire_430,
fourFunc_wire_431,
fourFunc_wire_432,
fourFunc_wire_433,
fourFunc_wire_434,
fourFunc_wire_435,
fourFunc_wire_436,
fourFunc_wire_437,
fourFunc_wire_438,
fourFunc_wire_439,
fourFunc_wire_440,
fourFunc_wire_441,
fourFunc_wire_442,
fourFunc_wire_443,
fourFunc_wire_444,
fourFunc_wire_445,
fourFunc_wire_446,
fourFunc_wire_447,
fourFunc_wire_448,
fourFunc_wire_449,
fourFunc_wire_450,
fourFunc_wire_451,
fourFunc_wire_452,
fourFunc_wire_453,
fourFunc_wire_454,
fourFunc_wire_455,
fourFunc_wire_456,
fourFunc_wire_457,
fourFunc_wire_458,
fourFunc_wire_459,
fourFunc_wire_460,
fourFunc_wire_461,
fourFunc_wire_462,
fourFunc_wire_463,
fourFunc_wire_464,
fourFunc_wire_465,
fourFunc_wire_466,
fourFunc_wire_467,
fourFunc_wire_468,
fourFunc_wire_469,
fourFunc_wire_470,
fourFunc_wire_471,
fourFunc_wire_472,
fourFunc_wire_473,
fourFunc_wire_474,
fourFunc_wire_475,
fourFunc_wire_476,
fourFunc_wire_477,
fourFunc_wire_478,
fourFunc_wire_479,
fourFunc_wire_480,
fourFunc_wire_481,
fourFunc_wire_482,
fourFunc_wire_483,
fourFunc_wire_484,
fourFunc_wire_485,
fourFunc_wire_486,
fourFunc_wire_487,
fourFunc_wire_488,
fourFunc_wire_489,
fourFunc_wire_490,
fourFunc_wire_491,
fourFunc_wire_492,
fourFunc_wire_493,
fourFunc_wire_494,
fourFunc_wire_495,
fourFunc_wire_496,
fourFunc_wire_497,
fourFunc_wire_498,
fourFunc_wire_499,
fourFunc_wire_500,
fourFunc_wire_501,
fourFunc_wire_502,
fourFunc_wire_503,
fourFunc_wire_504,
fourFunc_wire_505,
fourFunc_wire_506,
fourFunc_wire_507,
fourFunc_wire_508,
fourFunc_wire_509,
fourFunc_wire_510,
fourFunc_wire_511,
fourFunc_wire_512,
fourFunc_wire_513,
fourFunc_wire_514,
fourFunc_wire_515,
fourFunc_wire_516,
fourFunc_wire_517,
fourFunc_wire_518,
fourFunc_wire_519,
fourFunc_wire_520,
fourFunc_wire_521,
fourFunc_wire_522,
fourFunc_wire_523,
fourFunc_wire_524,
fourFunc_wire_525,
fourFunc_wire_526,
fourFunc_wire_527,
fourFunc_wire_528,
fourFunc_wire_529,
fourFunc_wire_530,
fourFunc_wire_531,
fourFunc_wire_532,
fourFunc_wire_533,
fourFunc_wire_534,
fourFunc_wire_535,
fourFunc_wire_536,
fourFunc_wire_537,
fourFunc_wire_538,
fourFunc_wire_539,
fourFunc_wire_540,
fourFunc_wire_541,
fourFunc_wire_542,
fourFunc_wire_543,
fourFunc_wire_544,
fourFunc_wire_545,
fourFunc_wire_546,
fourFunc_wire_547,
fourFunc_wire_548,
fourFunc_wire_549,
fourFunc_wire_550,
fourFunc_wire_551,
fourFunc_wire_552,
fourFunc_wire_553,
fourFunc_wire_554,
fourFunc_wire_555,
fourFunc_wire_556,
fourFunc_wire_557,
fourFunc_wire_558,
fourFunc_wire_559,
fourFunc_wire_560,
fourFunc_wire_561,
fourFunc_wire_562,
fourFunc_wire_563,
fourFunc_wire_564,
fourFunc_wire_565,
fourFunc_wire_566,
fourFunc_wire_567,
fourFunc_wire_568,
fourFunc_wire_569,
fourFunc_wire_570,
fourFunc_wire_571,
fourFunc_wire_572,
fourFunc_wire_573,
fourFunc_wire_574,
fourFunc_wire_575,
fourFunc_wire_576,
fourFunc_wire_577,
fourFunc_wire_578,
fourFunc_wire_579,
fourFunc_wire_580,
fourFunc_wire_581,
fourFunc_wire_582,
fourFunc_wire_583,
fourFunc_wire_584,
fourFunc_wire_585,
fourFunc_wire_586,
fourFunc_wire_587,
fourFunc_wire_588,
fourFunc_wire_589,
fourFunc_wire_590,
fourFunc_wire_591,
fourFunc_wire_592,
fourFunc_wire_593,
fourFunc_wire_594,
fourFunc_wire_595,
fourFunc_wire_596,
fourFunc_wire_597,
fourFunc_wire_598,
fourFunc_wire_599,
fourFunc_wire_600,
fourFunc_wire_601,
fourFunc_wire_602,
fourFunc_wire_603,
fourFunc_wire_604,
fourFunc_wire_605,
fourFunc_wire_606,
fourFunc_wire_607,
fourFunc_wire_608,
fourFunc_wire_609,
fourFunc_wire_610,
fourFunc_wire_611,
fourFunc_wire_612,
fourFunc_wire_613,
fourFunc_wire_614,
fourFunc_wire_615,
fourFunc_wire_616,
fourFunc_wire_617,
fourFunc_wire_618,
fourFunc_wire_619,
fourFunc_wire_620,
fourFunc_wire_621,
fourFunc_wire_622,
fourFunc_wire_623,
fourFunc_wire_624,
fourFunc_wire_625,
fourFunc_wire_626,
fourFunc_wire_627,
fourFunc_wire_628,
fourFunc_wire_629,
fourFunc_wire_630,
fourFunc_wire_631,
fourFunc_wire_632,
fourFunc_wire_633,
fourFunc_wire_634,
fourFunc_wire_635,
fourFunc_wire_636,
fourFunc_wire_637,
fourFunc_wire_638,
fourFunc_wire_639,
fourFunc_wire_640,
fourFunc_wire_641,
fourFunc_wire_642,
fourFunc_wire_643,
fourFunc_wire_644,
fourFunc_wire_645,
fourFunc_wire_646,
fourFunc_wire_647,
fourFunc_wire_648,
fourFunc_wire_649,
fourFunc_wire_650,
fourFunc_wire_651,
fourFunc_wire_652,
fourFunc_wire_653,
fourFunc_wire_654,
fourFunc_wire_655,
fourFunc_wire_656,
fourFunc_wire_657,
fourFunc_wire_658,
fourFunc_wire_659,
fourFunc_wire_660,
fourFunc_wire_661,
fourFunc_wire_662,
fourFunc_wire_663,
fourFunc_wire_664,
fourFunc_wire_665,
fourFunc_wire_666,
fourFunc_wire_667,
fourFunc_wire_668,
fourFunc_wire_669,
fourFunc_wire_670,
fourFunc_wire_671,
fourFunc_wire_672,
fourFunc_wire_673,
fourFunc_wire_674,
fourFunc_wire_675,
fourFunc_wire_676,
fourFunc_wire_677,
fourFunc_wire_678,
fourFunc_wire_679,
fourFunc_wire_680,
fourFunc_wire_681,
fourFunc_wire_682,
fourFunc_wire_683,
fourFunc_wire_684,
fourFunc_wire_685,
fourFunc_wire_686,
fourFunc_wire_687,
fourFunc_wire_688,
fourFunc_wire_689,
fourFunc_wire_690,
fourFunc_wire_691,
fourFunc_wire_692,
fourFunc_wire_693,
fourFunc_wire_694,
fourFunc_wire_695,
fourFunc_wire_696,
fourFunc_wire_697,
fourFunc_wire_698,
fourFunc_wire_699,
fourFunc_wire_700,
fourFunc_wire_701,
fourFunc_wire_702,
fourFunc_wire_703,
fourFunc_wire_704,
fourFunc_wire_705,
fourFunc_wire_706,
fourFunc_wire_707,
fourFunc_wire_708,
fourFunc_wire_709,
fourFunc_wire_710,
fourFunc_wire_711,
fourFunc_wire_712,
fourFunc_wire_713,
fourFunc_wire_714,
fourFunc_wire_715,
fourFunc_wire_716,
fourFunc_wire_717,
fourFunc_wire_718,
fourFunc_wire_719,
fourFunc_wire_720,
fourFunc_wire_721,
fourFunc_wire_722,
fourFunc_wire_723,
fourFunc_wire_724,
fourFunc_wire_725,
fourFunc_wire_726,
fourFunc_wire_727,
fourFunc_wire_728,
fourFunc_wire_729,
fourFunc_wire_730,
fourFunc_wire_731,
fourFunc_wire_732,
fourFunc_wire_733,
fourFunc_wire_734,
fourFunc_wire_735,
fourFunc_wire_736,
fourFunc_wire_737,
fourFunc_wire_738,
fourFunc_wire_739,
fourFunc_wire_740,
fourFunc_wire_741,
fourFunc_wire_742,
fourFunc_wire_743,
fourFunc_wire_744,
fourFunc_wire_745,
fourFunc_wire_746,
fourFunc_wire_747,
fourFunc_wire_748,
fourFunc_wire_749,
fourFunc_wire_750,
fourFunc_wire_751,
fourFunc_wire_752,
fourFunc_wire_753,
fourFunc_wire_754,
fourFunc_wire_755,
fourFunc_wire_756,
fourFunc_wire_757,
fourFunc_wire_758,
fourFunc_wire_759,
fourFunc_wire_760,
fourFunc_wire_761,
fourFunc_wire_762,
fourFunc_wire_763,
fourFunc_wire_764,
fourFunc_wire_765,
fourFunc_wire_766,
fourFunc_wire_767,
fourFunc_wire_768,
fourFunc_wire_769,
fourFunc_wire_770,
fourFunc_wire_771,
fourFunc_wire_772,
fourFunc_wire_773,
fourFunc_wire_774,
fourFunc_wire_775,
fourFunc_wire_776,
fourFunc_wire_777,
fourFunc_wire_778,
fourFunc_wire_779,
fourFunc_wire_780,
fourFunc_wire_781,
fourFunc_wire_782,
fourFunc_wire_783,
fourFunc_wire_784,
fourFunc_wire_785,
fourFunc_wire_786,
fourFunc_wire_787,
fourFunc_wire_788,
fourFunc_wire_789,
fourFunc_wire_790,
fourFunc_wire_791,
fourFunc_wire_792,
fourFunc_wire_793,
fourFunc_wire_794,
fourFunc_wire_795,
fourFunc_wire_796,
fourFunc_wire_797,
fourFunc_wire_798,
fourFunc_wire_799,
fourFunc_wire_800,
fourFunc_wire_801,
fourFunc_wire_802,
fourFunc_wire_803,
fourFunc_wire_804,
fourFunc_wire_805,
fourFunc_wire_806,
fourFunc_wire_807,
fourFunc_wire_808,
fourFunc_wire_809,
fourFunc_wire_810,
fourFunc_wire_811,
fourFunc_wire_812,
fourFunc_wire_813,
fourFunc_wire_814,
fourFunc_wire_815,
fourFunc_wire_816,
fourFunc_wire_817,
fourFunc_wire_818,
fourFunc_wire_819,
fourFunc_wire_820,
fourFunc_wire_821,
fourFunc_wire_822,
fourFunc_wire_823,
fourFunc_wire_824,
fourFunc_wire_825,
fourFunc_wire_826,
fourFunc_wire_827,
fourFunc_wire_828,
fourFunc_wire_829,
fourFunc_wire_830,
fourFunc_wire_831,
fourFunc_wire_832,
fourFunc_wire_833,
fourFunc_wire_834,
fourFunc_wire_835,
fourFunc_wire_836,
fourFunc_wire_837,
fourFunc_wire_838,
fourFunc_wire_839,
fourFunc_wire_840,
fourFunc_wire_841,
fourFunc_wire_842,
fourFunc_wire_843,
fourFunc_wire_844,
fourFunc_wire_845,
fourFunc_wire_846,
fourFunc_wire_847,
fourFunc_wire_848,
fourFunc_wire_849,
fourFunc_wire_850,
fourFunc_wire_851,
fourFunc_wire_852,
fourFunc_wire_853,
fourFunc_wire_854,
fourFunc_wire_855,
fourFunc_wire_856,
fourFunc_wire_857,
fourFunc_wire_858,
fourFunc_wire_35_0,
fourFunc_wire_35_1,
fourFunc_wire_46_0,
fourFunc_wire_46_1,
fourFunc_wire_122_0,
fourFunc_wire_122_1,
fourFunc_wire_122_2,
fourFunc_wire_133_0,
fourFunc_wire_133_1,
fourFunc_wire_133_2,
fourFunc_wire_138_0,
fourFunc_wire_138_1,
fourFunc_wire_138_2,
fourFunc_wire_143_0,
fourFunc_wire_143_1,
fourFunc_wire_143_2,
fourFunc_wire_148_0,
fourFunc_wire_148_1,
fourFunc_wire_148_2,
fourFunc_wire_153_0,
fourFunc_wire_153_1,
fourFunc_wire_153_2,
fourFunc_wire_158_0,
fourFunc_wire_158_1,
fourFunc_wire_158_2,
fourFunc_wire_184_0,
fourFunc_wire_184_1,
fourFunc_wire_166_0,
fourFunc_wire_166_1,
fourFunc_wire_166_2,
fourFunc_wire_170_0,
fourFunc_wire_170_1,
fourFunc_wire_170_2,
fourFunc_wire_174_0,
fourFunc_wire_174_1,
fourFunc_wire_174_2,
fourFunc_wire_178_0,
fourFunc_wire_178_1,
fourFunc_wire_178_2,
fourFunc_wire_182_0,
fourFunc_wire_182_1,
fourFunc_wire_182_2,
fourFunc_wire_187_0,
fourFunc_wire_187_1,
fourFunc_wire_187_2,
fourFunc_wire_213_0,
fourFunc_wire_213_1,
fourFunc_wire_195_0,
fourFunc_wire_195_1,
fourFunc_wire_195_2,
fourFunc_wire_199_0,
fourFunc_wire_199_1,
fourFunc_wire_199_2,
fourFunc_wire_203_0,
fourFunc_wire_203_1,
fourFunc_wire_203_2,
fourFunc_wire_207_0,
fourFunc_wire_207_1,
fourFunc_wire_207_2,
fourFunc_wire_211_0,
fourFunc_wire_211_1,
fourFunc_wire_211_2,
fourFunc_wire_216_0,
fourFunc_wire_216_1,
fourFunc_wire_216_2,
fourFunc_wire_242_0,
fourFunc_wire_242_1,
fourFunc_wire_224_0,
fourFunc_wire_224_1,
fourFunc_wire_224_2,
fourFunc_wire_228_0,
fourFunc_wire_228_1,
fourFunc_wire_228_2,
fourFunc_wire_232_0,
fourFunc_wire_232_1,
fourFunc_wire_232_2,
fourFunc_wire_236_0,
fourFunc_wire_236_1,
fourFunc_wire_236_2,
fourFunc_wire_240_0,
fourFunc_wire_240_1,
fourFunc_wire_240_2,
fourFunc_wire_245_0,
fourFunc_wire_245_1,
fourFunc_wire_245_2,
fourFunc_wire_271_0,
fourFunc_wire_271_1,
fourFunc_wire_253_0,
fourFunc_wire_253_1,
fourFunc_wire_253_2,
fourFunc_wire_257_0,
fourFunc_wire_257_1,
fourFunc_wire_257_2,
fourFunc_wire_261_0,
fourFunc_wire_261_1,
fourFunc_wire_261_2,
fourFunc_wire_265_0,
fourFunc_wire_265_1,
fourFunc_wire_265_2,
fourFunc_wire_269_0,
fourFunc_wire_269_1,
fourFunc_wire_269_2,
fourFunc_wire_274_0,
fourFunc_wire_274_1,
fourFunc_wire_274_2,
fourFunc_wire_299_0,
fourFunc_wire_299_1,
fourFunc_wire_285_0,
fourFunc_wire_285_1,
fourFunc_wire_285_2,
fourFunc_wire_289_0,
fourFunc_wire_289_1,
fourFunc_wire_289_2,
fourFunc_wire_293_0,
fourFunc_wire_293_1,
fourFunc_wire_293_2,
fourFunc_wire_297_0,
fourFunc_wire_297_1,
fourFunc_wire_297_2,
fourFunc_wire_302_0,
fourFunc_wire_302_1,
fourFunc_wire_302_2,
fourFunc_wire_324_0,
fourFunc_wire_324_1,
fourFunc_wire_121_0,
fourFunc_wire_121_1,
fourFunc_wire_118_0,
fourFunc_wire_118_1,
fourFunc_wire_115_0,
fourFunc_wire_115_1,
fourFunc_wire_112_0,
fourFunc_wire_112_1,
fourFunc_wire_109_0,
fourFunc_wire_109_1,
fourFunc_wire_106_0,
fourFunc_wire_106_1,
fourFunc_wire_103_0,
fourFunc_wire_103_1,
fourFunc_wire_98_0,
fourFunc_wire_98_1,
fourFunc_wire_306_0,
fourFunc_wire_306_1,
fourFunc_wire_310_0,
fourFunc_wire_310_1,
fourFunc_wire_314_0,
fourFunc_wire_314_1,
fourFunc_wire_318_0,
fourFunc_wire_318_1,
fourFunc_wire_322_0,
fourFunc_wire_322_1,
fourFunc_wire_327_0,
fourFunc_wire_327_1,
fourFunc_wire_278_0,
fourFunc_wire_278_1,
fourFunc_wire_278_2,
fourFunc_wire_124_0,
fourFunc_wire_124_1,
fourFunc_wire_307_0,
fourFunc_wire_307_1,
fourFunc_wire_307_2,
fourFunc_wire_311_0,
fourFunc_wire_311_1,
fourFunc_wire_311_2,
fourFunc_wire_315_0,
fourFunc_wire_315_1,
fourFunc_wire_315_2,
fourFunc_wire_319_0,
fourFunc_wire_319_1,
fourFunc_wire_319_2,
fourFunc_wire_323_0,
fourFunc_wire_323_1,
fourFunc_wire_323_2,
fourFunc_wire_328_0,
fourFunc_wire_328_1,
fourFunc_wire_279_0,
fourFunc_wire_279_1,
fourFunc_wire_282_0,
fourFunc_wire_282_1,
fourFunc_wire_286_0,
fourFunc_wire_286_1,
fourFunc_wire_290_0,
fourFunc_wire_290_1,
fourFunc_wire_294_0,
fourFunc_wire_294_1,
fourFunc_wire_298_0,
fourFunc_wire_298_1,
fourFunc_wire_250_0,
fourFunc_wire_250_1,
fourFunc_wire_254_0,
fourFunc_wire_254_1,
fourFunc_wire_258_0,
fourFunc_wire_258_1,
fourFunc_wire_262_0,
fourFunc_wire_262_1,
fourFunc_wire_266_0,
fourFunc_wire_266_1,
fourFunc_wire_270_0,
fourFunc_wire_270_1,
fourFunc_wire_221_0,
fourFunc_wire_221_1,
fourFunc_wire_225_0,
fourFunc_wire_225_1,
fourFunc_wire_229_0,
fourFunc_wire_229_1,
fourFunc_wire_233_0,
fourFunc_wire_233_1,
fourFunc_wire_237_0,
fourFunc_wire_237_1,
fourFunc_wire_241_0,
fourFunc_wire_241_1,
fourFunc_wire_192_0,
fourFunc_wire_192_1,
fourFunc_wire_196_0,
fourFunc_wire_196_1,
fourFunc_wire_200_0,
fourFunc_wire_200_1,
fourFunc_wire_204_0,
fourFunc_wire_204_1,
fourFunc_wire_208_0,
fourFunc_wire_208_1,
fourFunc_wire_212_0,
fourFunc_wire_212_1,
fourFunc_wire_163_0,
fourFunc_wire_163_1,
fourFunc_wire_167_0,
fourFunc_wire_167_1,
fourFunc_wire_171_0,
fourFunc_wire_171_1,
fourFunc_wire_175_0,
fourFunc_wire_175_1,
fourFunc_wire_179_0,
fourFunc_wire_179_1,
fourFunc_wire_183_0,
fourFunc_wire_183_1,
fourFunc_wire_129_0,
fourFunc_wire_129_1,
fourFunc_wire_134_0,
fourFunc_wire_134_1,
fourFunc_wire_139_0,
fourFunc_wire_139_1,
fourFunc_wire_144_0,
fourFunc_wire_144_1,
fourFunc_wire_149_0,
fourFunc_wire_149_1,
fourFunc_wire_154_0,
fourFunc_wire_154_1,
fourFunc_wire_249_0,
fourFunc_wire_249_1,
fourFunc_wire_249_2,
fourFunc_wire_220_0,
fourFunc_wire_220_1,
fourFunc_wire_220_2,
fourFunc_wire_191_0,
fourFunc_wire_191_1,
fourFunc_wire_191_2,
fourFunc_wire_162_0,
fourFunc_wire_162_1,
fourFunc_wire_162_2,
fourFunc_wire_128_0,
fourFunc_wire_128_1,
fourFunc_wire_128_2,
fourFunc_wire_321_0,
fourFunc_wire_321_1,
fourFunc_wire_321_2,
fourFunc_wire_317_0,
fourFunc_wire_317_1,
fourFunc_wire_317_2,
fourFunc_wire_313_0,
fourFunc_wire_313_1,
fourFunc_wire_313_2,
fourFunc_wire_309_0,
fourFunc_wire_309_1,
fourFunc_wire_309_2,
fourFunc_wire_305_0,
fourFunc_wire_305_1,
fourFunc_wire_305_2,
fourFunc_wire_123_0,
fourFunc_wire_123_1,
fourFunc_wire_296_0,
fourFunc_wire_296_1,
fourFunc_wire_296_2,
fourFunc_wire_292_0,
fourFunc_wire_292_1,
fourFunc_wire_292_2,
fourFunc_wire_288_0,
fourFunc_wire_288_1,
fourFunc_wire_288_2,
fourFunc_wire_284_0,
fourFunc_wire_284_1,
fourFunc_wire_284_2,
fourFunc_wire_281_0,
fourFunc_wire_281_1,
fourFunc_wire_281_2,
fourFunc_wire_277_0,
fourFunc_wire_277_1,
fourFunc_wire_277_2,
fourFunc_wire_268_0,
fourFunc_wire_268_1,
fourFunc_wire_268_2,
fourFunc_wire_264_0,
fourFunc_wire_264_1,
fourFunc_wire_264_2,
fourFunc_wire_260_0,
fourFunc_wire_260_1,
fourFunc_wire_260_2,
fourFunc_wire_256_0,
fourFunc_wire_256_1,
fourFunc_wire_256_2,
fourFunc_wire_252_0,
fourFunc_wire_252_1,
fourFunc_wire_252_2,
fourFunc_wire_248_0,
fourFunc_wire_248_1,
fourFunc_wire_248_2,
fourFunc_wire_239_0,
fourFunc_wire_239_1,
fourFunc_wire_239_2,
fourFunc_wire_235_0,
fourFunc_wire_235_1,
fourFunc_wire_235_2,
fourFunc_wire_231_0,
fourFunc_wire_231_1,
fourFunc_wire_231_2,
fourFunc_wire_227_0,
fourFunc_wire_227_1,
fourFunc_wire_227_2,
fourFunc_wire_223_0,
fourFunc_wire_223_1,
fourFunc_wire_223_2,
fourFunc_wire_219_0,
fourFunc_wire_219_1,
fourFunc_wire_219_2,
fourFunc_wire_210_0,
fourFunc_wire_210_1,
fourFunc_wire_210_2,
fourFunc_wire_206_0,
fourFunc_wire_206_1,
fourFunc_wire_206_2,
fourFunc_wire_202_0,
fourFunc_wire_202_1,
fourFunc_wire_202_2,
fourFunc_wire_198_0,
fourFunc_wire_198_1,
fourFunc_wire_198_2,
fourFunc_wire_194_0,
fourFunc_wire_194_1,
fourFunc_wire_194_2,
fourFunc_wire_190_0,
fourFunc_wire_190_1,
fourFunc_wire_190_2,
fourFunc_wire_181_0,
fourFunc_wire_181_1,
fourFunc_wire_181_2,
fourFunc_wire_177_0,
fourFunc_wire_177_1,
fourFunc_wire_177_2,
fourFunc_wire_173_0,
fourFunc_wire_173_1,
fourFunc_wire_173_2,
fourFunc_wire_169_0,
fourFunc_wire_169_1,
fourFunc_wire_169_2,
fourFunc_wire_165_0,
fourFunc_wire_165_1,
fourFunc_wire_165_2,
fourFunc_wire_161_0,
fourFunc_wire_161_1,
fourFunc_wire_161_2,
fourFunc_wire_152_0,
fourFunc_wire_152_1,
fourFunc_wire_152_2,
fourFunc_wire_147_0,
fourFunc_wire_147_1,
fourFunc_wire_147_2,
fourFunc_wire_142_0,
fourFunc_wire_142_1,
fourFunc_wire_142_2,
fourFunc_wire_137_0,
fourFunc_wire_137_1,
fourFunc_wire_137_2,
fourFunc_wire_132_0,
fourFunc_wire_132_1,
fourFunc_wire_132_2,
fourFunc_wire_127_0,
fourFunc_wire_127_1,
fourFunc_wire_127_2,
fourFunc_wire_93_0,
fourFunc_wire_93_1,
fourFunc_wire_88_0,
fourFunc_wire_88_1,
fourFunc_wire_83_0,
fourFunc_wire_83_1,
fourFunc_wire_78_0,
fourFunc_wire_78_1,
fourFunc_wire_73_0,
fourFunc_wire_73_1,
fourFunc_wire_68_0,
fourFunc_wire_68_1,
fourFunc_wire_63_0,
fourFunc_wire_63_1,
fourFunc_wire_60_0,
fourFunc_wire_60_1,
fourFunc_wire_551_0,
fourFunc_wire_551_1,
fourFunc_wire_551_2,
fourFunc_wire_551_3,
fourFunc_wire_551_4,
fourFunc_wire_551_5,
fourFunc_wire_551_6,
fourFunc_wire_551_7,
fourFunc_wire_551_8,
fourFunc_wire_551_9,
fourFunc_wire_551_10,
fourFunc_wire_551_11,
fourFunc_wire_551_12,
fourFunc_wire_551_13,
fourFunc_wire_551_14,
fourFunc_wire_551_15,
fourFunc_wire_551_16,
fourFunc_wire_551_17,
fourFunc_wire_551_18,
fourFunc_wire_551_19,
fourFunc_wire_551_20,
fourFunc_wire_551_21,
fourFunc_wire_2_0,
fourFunc_wire_2_1,
fourFunc_wire_2_2,
fourFunc_wire_2_3,
fourFunc_wire_2_4,
fourFunc_wire_2_5,
fourFunc_wire_2_6,
fourFunc_wire_2_7,
fourFunc_wire_2_8,
fourFunc_wire_2_9,
fourFunc_wire_2_10,
fourFunc_wire_10_0,
fourFunc_wire_10_1,
fourFunc_wire_10_2,
fourFunc_wire_10_3,
fourFunc_wire_10_4,
fourFunc_wire_10_5,
fourFunc_wire_10_6,
fourFunc_wire_10_7,
fourFunc_wire_10_8,
fourFunc_wire_10_9,
fourFunc_wire_10_10,
fourFunc_wire_3_0,
fourFunc_wire_3_1,
fourFunc_wire_3_2,
fourFunc_wire_3_3,
fourFunc_wire_3_4,
fourFunc_wire_3_5,
fourFunc_wire_3_6,
fourFunc_wire_3_7,
fourFunc_wire_3_8,
fourFunc_wire_8_0,
fourFunc_wire_8_1,
fourFunc_wire_8_2,
fourFunc_wire_8_3,
fourFunc_wire_8_4,
fourFunc_wire_8_5,
fourFunc_wire_8_6,
fourFunc_wire_8_7,
fourFunc_wire_8_8,
fourFunc_wire_8_9,
fourFunc_wire_8_10,
fourFunc_wire_8_11,
fourFunc_wire_552_0,
fourFunc_wire_552_1,
fourFunc_wire_553_0,
fourFunc_wire_553_1,
fourFunc_wire_554_0,
fourFunc_wire_554_1,
fourFunc_wire_555_0,
fourFunc_wire_555_1,
fourFunc_wire_556_0,
fourFunc_wire_556_1,
fourFunc_wire_557_0,
fourFunc_wire_557_1,
fourFunc_wire_558_0,
fourFunc_wire_558_1,
fourFunc_wire_559_0,
fourFunc_wire_559_1,
fourFunc_wire_53_0,
fourFunc_wire_53_1,
fourFunc_wire_53_2,
fourFunc_wire_53_3,
fourFunc_wire_53_4,
fourFunc_wire_53_5,
fourFunc_wire_53_6,
fourFunc_wire_53_7,
fourFunc_wire_53_8,
fourFunc_wire_53_9,
fourFunc_wire_53_10,
fourFunc_wire_53_11,
fourFunc_wire_53_12,
fourFunc_wire_53_13,
fourFunc_wire_53_14,
fourFunc_wire_53_15,
fourFunc_wire_53_16,
fourFunc_wire_53_17,
fourFunc_wire_53_18,
fourFunc_wire_95_0,
fourFunc_wire_95_1,
fourFunc_wire_95_2,
fourFunc_wire_95_3,
fourFunc_wire_95_4,
fourFunc_wire_95_5,
fourFunc_wire_95_6,
fourFunc_wire_95_7,
fourFunc_wire_95_8,
fourFunc_wire_95_9,
fourFunc_wire_95_10,
fourFunc_wire_95_11,
fourFunc_wire_95_12,
fourFunc_wire_95_13,
fourFunc_wire_95_14,
fourFunc_wire_95_15,
fourFunc_wire_95_16,
fourFunc_wire_95_17,
fourFunc_wire_95_18,
fourFunc_wire_95_19,
fourFunc_wire_95_20,
fourFunc_wire_95_21,
fourFunc_wire_95_22,
fourFunc_wire_95_23,
fourFunc_wire_95_24,
fourFunc_wire_95_25,
fourFunc_wire_95_26,
fourFunc_wire_95_27,
fourFunc_wire_90_0,
fourFunc_wire_90_1,
fourFunc_wire_90_2,
fourFunc_wire_90_3,
fourFunc_wire_90_4,
fourFunc_wire_90_5,
fourFunc_wire_90_6,
fourFunc_wire_90_7,
fourFunc_wire_90_8,
fourFunc_wire_90_9,
fourFunc_wire_90_10,
fourFunc_wire_90_11,
fourFunc_wire_90_12,
fourFunc_wire_90_13,
fourFunc_wire_90_14,
fourFunc_wire_85_0,
fourFunc_wire_85_1,
fourFunc_wire_85_2,
fourFunc_wire_85_3,
fourFunc_wire_85_4,
fourFunc_wire_85_5,
fourFunc_wire_85_6,
fourFunc_wire_85_7,
fourFunc_wire_85_8,
fourFunc_wire_85_9,
fourFunc_wire_85_10,
fourFunc_wire_85_11,
fourFunc_wire_85_12,
fourFunc_wire_85_13,
fourFunc_wire_85_14,
fourFunc_wire_80_0,
fourFunc_wire_80_1,
fourFunc_wire_80_2,
fourFunc_wire_80_3,
fourFunc_wire_80_4,
fourFunc_wire_80_5,
fourFunc_wire_80_6,
fourFunc_wire_80_7,
fourFunc_wire_80_8,
fourFunc_wire_80_9,
fourFunc_wire_80_10,
fourFunc_wire_80_11,
fourFunc_wire_80_12,
fourFunc_wire_80_13,
fourFunc_wire_80_14,
fourFunc_wire_75_0,
fourFunc_wire_75_1,
fourFunc_wire_75_2,
fourFunc_wire_75_3,
fourFunc_wire_75_4,
fourFunc_wire_75_5,
fourFunc_wire_75_6,
fourFunc_wire_75_7,
fourFunc_wire_75_8,
fourFunc_wire_75_9,
fourFunc_wire_75_10,
fourFunc_wire_75_11,
fourFunc_wire_75_12,
fourFunc_wire_75_13,
fourFunc_wire_75_14,
fourFunc_wire_70_0,
fourFunc_wire_70_1,
fourFunc_wire_70_2,
fourFunc_wire_70_3,
fourFunc_wire_70_4,
fourFunc_wire_70_5,
fourFunc_wire_70_6,
fourFunc_wire_70_7,
fourFunc_wire_70_8,
fourFunc_wire_70_9,
fourFunc_wire_70_10,
fourFunc_wire_70_11,
fourFunc_wire_70_12,
fourFunc_wire_70_13,
fourFunc_wire_70_14,
fourFunc_wire_65_0,
fourFunc_wire_65_1,
fourFunc_wire_65_2,
fourFunc_wire_65_3,
fourFunc_wire_65_4,
fourFunc_wire_65_5,
fourFunc_wire_65_6,
fourFunc_wire_65_7,
fourFunc_wire_65_8,
fourFunc_wire_65_9,
fourFunc_wire_65_10,
fourFunc_wire_65_11,
fourFunc_wire_65_12,
fourFunc_wire_65_13,
fourFunc_wire_65_14,
fourFunc_wire_54_0,
fourFunc_wire_54_1,
fourFunc_wire_54_2,
fourFunc_wire_54_3,
fourFunc_wire_54_4,
fourFunc_wire_54_5,
fourFunc_wire_94_0,
fourFunc_wire_94_1,
fourFunc_wire_94_2,
fourFunc_wire_94_3,
fourFunc_wire_94_4,
fourFunc_wire_94_5,
fourFunc_wire_94_6,
fourFunc_wire_94_7,
fourFunc_wire_89_0,
fourFunc_wire_89_1,
fourFunc_wire_89_2,
fourFunc_wire_89_3,
fourFunc_wire_89_4,
fourFunc_wire_89_5,
fourFunc_wire_89_6,
fourFunc_wire_89_7,
fourFunc_wire_84_0,
fourFunc_wire_84_1,
fourFunc_wire_84_2,
fourFunc_wire_84_3,
fourFunc_wire_84_4,
fourFunc_wire_84_5,
fourFunc_wire_84_6,
fourFunc_wire_84_7,
fourFunc_wire_79_0,
fourFunc_wire_79_1,
fourFunc_wire_79_2,
fourFunc_wire_79_3,
fourFunc_wire_79_4,
fourFunc_wire_79_5,
fourFunc_wire_79_6,
fourFunc_wire_79_7,
fourFunc_wire_74_0,
fourFunc_wire_74_1,
fourFunc_wire_74_2,
fourFunc_wire_74_3,
fourFunc_wire_74_4,
fourFunc_wire_74_5,
fourFunc_wire_74_6,
fourFunc_wire_74_7,
fourFunc_wire_69_0,
fourFunc_wire_69_1,
fourFunc_wire_69_2,
fourFunc_wire_69_3,
fourFunc_wire_69_4,
fourFunc_wire_69_5,
fourFunc_wire_69_6,
fourFunc_wire_69_7,
fourFunc_wire_64_0,
fourFunc_wire_64_1,
fourFunc_wire_64_2,
fourFunc_wire_64_3,
fourFunc_wire_64_4,
fourFunc_wire_64_5,
fourFunc_wire_64_6,
fourFunc_wire_64_7,
fourFunc_wire_59_0,
fourFunc_wire_59_1,
fourFunc_wire_59_2,
fourFunc_wire_59_3,
fourFunc_wire_59_4,
fourFunc_wire_59_5,
fourFunc_wire_56_0,
fourFunc_wire_56_1,
fourFunc_wire_56_2,
fourFunc_wire_56_3,
fourFunc_wire_582_0,
fourFunc_wire_582_1,
fourFunc_wire_588_0,
fourFunc_wire_588_1,
fourFunc_wire_588_2,
fourFunc_wire_588_3,
fourFunc_wire_589_0,
fourFunc_wire_589_1,
fourFunc_wire_589_2,
fourFunc_wire_589_3,
fourFunc_wire_589_4,
fourFunc_wire_590_0,
fourFunc_wire_590_1,
fourFunc_wire_590_2,
fourFunc_wire_586_0,
fourFunc_wire_586_1,
fourFunc_wire_586_2,
fourFunc_wire_586_3,
fourFunc_wire_586_4,
fourFunc_wire_586_5,
fourFunc_wire_586_6,
fourFunc_wire_586_7,
fourFunc_wire_586_8,
fourFunc_wire_586_9,
fourFunc_wire_586_10,
fourFunc_wire_586_11,
fourFunc_wire_586_12,
fourFunc_wire_586_13,
fourFunc_wire_586_14,
fourFunc_wire_586_15,
fourFunc_wire_586_16,
fourFunc_wire_586_17,
fourFunc_wire_581_0,
fourFunc_wire_581_1,
fourFunc_wire_581_2,
fourFunc_wire_581_3,
fourFunc_wire_581_4,
fourFunc_wire_599_0,
fourFunc_wire_599_1,
fourFunc_wire_599_2,
fourFunc_wire_599_3,
fourFunc_wire_599_4,
fourFunc_wire_599_5,
fourFunc_wire_599_6,
fourFunc_wire_599_7,
fourFunc_wire_599_8,
fourFunc_wire_599_9,
fourFunc_wire_599_10,
fourFunc_wire_599_11,
fourFunc_wire_599_12,
fourFunc_wire_599_13,
fourFunc_wire_599_14,
fourFunc_wire_599_15,
fourFunc_wire_599_16,
fourFunc_wire_599_17,
fourFunc_wire_599_18,
fourFunc_wire_599_19,
fourFunc_wire_599_20,
fourFunc_wire_599_21,
fourFunc_wire_599_22,
fourFunc_wire_599_23,
fourFunc_wire_599_24,
fourFunc_wire_599_25,
fourFunc_wire_599_26,
fourFunc_wire_599_27,
fourFunc_wire_599_28,
fourFunc_wire_599_29,
fourFunc_wire_599_30,
fourFunc_wire_599_31,
fourFunc_wire_50_0,
fourFunc_wire_50_1,
fourFunc_wire_605_0,
fourFunc_wire_605_1,
fourFunc_wire_609_0,
fourFunc_wire_609_1,
fourFunc_wire_609_2,
fourFunc_wire_609_3,
fourFunc_wire_608_0,
fourFunc_wire_608_1,
fourFunc_wire_608_2,
fourFunc_wire_608_3,
fourFunc_wire_608_4,
fourFunc_wire_608_5,
fourFunc_wire_608_6,
fourFunc_wire_608_7,
fourFunc_wire_608_8,
fourFunc_wire_608_9,
fourFunc_wire_608_10,
fourFunc_wire_608_11,
fourFunc_wire_608_12,
fourFunc_wire_604_0,
fourFunc_wire_604_1,
fourFunc_wire_604_2,
fourFunc_wire_604_3,
fourFunc_wire_604_4,
fourFunc_wire_604_5,
fourFunc_wire_604_6,
fourFunc_wire_604_7,
fourFunc_wire_604_8,
fourFunc_wire_604_9,
fourFunc_wire_604_10,
fourFunc_wire_604_11,
fourFunc_wire_604_12,
fourFunc_wire_604_13,
fourFunc_wire_604_14,
fourFunc_wire_604_15,
fourFunc_wire_604_16,
fourFunc_wire_604_17,
fourFunc_wire_604_18,
fourFunc_wire_604_19,
fourFunc_wire_604_20,
fourFunc_wire_604_21,
fourFunc_wire_604_22,
fourFunc_wire_604_23,
fourFunc_wire_604_24,
fourFunc_wire_604_25,
fourFunc_wire_604_26,
fourFunc_wire_604_27,
fourFunc_wire_604_28,
fourFunc_wire_604_29,
fourFunc_wire_604_30,
fourFunc_wire_604_31,
fourFunc_wire_604_32,
fourFunc_wire_604_33,
fourFunc_wire_604_34,
fourFunc_wire_604_35,
fourFunc_wire_604_36,
fourFunc_wire_604_37,
fourFunc_wire_604_38,
fourFunc_wire_604_39,
fourFunc_wire_648_0,
fourFunc_wire_648_1,
fourFunc_wire_648_2,
fourFunc_wire_648_3,
fourFunc_wire_648_4,
fourFunc_wire_648_5,
fourFunc_wire_648_6,
fourFunc_wire_648_7,
fourFunc_wire_648_8,
fourFunc_wire_648_9,
fourFunc_wire_648_10,
fourFunc_wire_434_0,
fourFunc_wire_434_1,
fourFunc_wire_434_2,
fourFunc_wire_434_3,
fourFunc_wire_434_4,
fourFunc_wire_434_5,
fourFunc_wire_434_6,
fourFunc_wire_434_7,
fourFunc_wire_446_0,
fourFunc_wire_446_1,
fourFunc_wire_446_2,
fourFunc_wire_446_3,
fourFunc_wire_446_4,
fourFunc_wire_446_5,
fourFunc_wire_446_6,
fourFunc_wire_446_7,
fourFunc_wire_446_8,
fourFunc_wire_350_0,
fourFunc_wire_350_1,
fourFunc_wire_350_2,
fourFunc_wire_350_3,
fourFunc_wire_350_4,
fourFunc_wire_350_5,
fourFunc_wire_350_6,
fourFunc_wire_350_7,
fourFunc_wire_350_8,
fourFunc_wire_364_0,
fourFunc_wire_364_1,
fourFunc_wire_364_2,
fourFunc_wire_364_3,
fourFunc_wire_364_4,
fourFunc_wire_364_5,
fourFunc_wire_364_6,
fourFunc_wire_364_7,
fourFunc_wire_364_8,
fourFunc_wire_378_0,
fourFunc_wire_378_1,
fourFunc_wire_378_2,
fourFunc_wire_378_3,
fourFunc_wire_378_4,
fourFunc_wire_378_5,
fourFunc_wire_378_6,
fourFunc_wire_378_7,
fourFunc_wire_378_8,
fourFunc_wire_392_0,
fourFunc_wire_392_1,
fourFunc_wire_392_2,
fourFunc_wire_392_3,
fourFunc_wire_392_4,
fourFunc_wire_392_5,
fourFunc_wire_392_6,
fourFunc_wire_392_7,
fourFunc_wire_392_8,
fourFunc_wire_406_0,
fourFunc_wire_406_1,
fourFunc_wire_406_2,
fourFunc_wire_406_3,
fourFunc_wire_406_4,
fourFunc_wire_406_5,
fourFunc_wire_406_6,
fourFunc_wire_406_7,
fourFunc_wire_406_8,
fourFunc_wire_420_0,
fourFunc_wire_420_1,
fourFunc_wire_420_2,
fourFunc_wire_420_3,
fourFunc_wire_420_4,
fourFunc_wire_420_5,
fourFunc_wire_420_6,
fourFunc_wire_420_7,
fourFunc_wire_420_8,
fourFunc_wire_717_0,
fourFunc_wire_717_1,
fourFunc_wire_717_2,
fourFunc_wire_717_3,
fourFunc_wire_717_4,
fourFunc_wire_717_5,
fourFunc_wire_717_6,
fourFunc_wire_717_7,
fourFunc_wire_717_8,
fourFunc_wire_9_0,
fourFunc_wire_9_1,
fourFunc_wire_9_2,
fourFunc_wire_9_3,
fourFunc_wire_9_4,
fourFunc_wire_9_5,
fourFunc_wire_9_6,
fourFunc_wire_9_7,
fourFunc_wire_9_8,
fourFunc_wire_9_9,
fourFunc_wire_9_10,
fourFunc_wire_9_11,
fourFunc_wire_9_12,
fourFunc_wire_9_13,
fourFunc_wire_9_14,
fourFunc_wire_9_15,
fourFunc_wire_9_16,
fourFunc_wire_9_17,
fourFunc_wire_9_18,
fourFunc_wire_9_19,
fourFunc_wire_9_20,
fourFunc_wire_9_21,
fourFunc_wire_9_22,
fourFunc_wire_9_23,
fourFunc_wire_598_0,
fourFunc_wire_598_1,
fourFunc_wire_598_2,
fourFunc_wire_598_3,
fourFunc_wire_598_4,
fourFunc_wire_598_5,
fourFunc_wire_641_0,
fourFunc_wire_641_1,
fourFunc_wire_641_2,
fourFunc_wire_626_0,
fourFunc_wire_626_1,
fourFunc_wire_626_2,
fourFunc_wire_628_0,
fourFunc_wire_628_1,
fourFunc_wire_628_2,
fourFunc_wire_630_0,
fourFunc_wire_630_1,
fourFunc_wire_630_2,
fourFunc_wire_634_0,
fourFunc_wire_634_1,
fourFunc_wire_634_2,
fourFunc_wire_636_0,
fourFunc_wire_636_1,
fourFunc_wire_636_2,
fourFunc_wire_632_0,
fourFunc_wire_632_1,
fourFunc_wire_632_2,
fourFunc_wire_638_0,
fourFunc_wire_638_1,
fourFunc_wire_638_2,
fourFunc_wire_640_0,
fourFunc_wire_640_1,
fourFunc_wire_640_2,
NOT_intermediateXXXwire_690_0,
NOT_intermediateXXXwire_690_1,
NOT_intermediateXXXwire_690_2,
NOT_intermediateXXXwire_697_0,
NOT_intermediateXXXwire_697_1,
NOT_intermediateXXXwire_697_2,
NOT_intermediateXXXwire_697_3,
NOT_intermediateXXXwire_697_4,
NOT_intermediateXXXwire_697_5,
NOT_intermediateXXXwire_697_6,
NOT_intermediateXXXwire_697_7,
NOT_intermediateXXXwire_922_0,
NOT_intermediateXXXwire_922_1,
NOT_intermediateXXXwire_922_2,
NOT_intermediateXXXwire_922_3,
NOT_intermediateXXXwire_922_4,
NOT_intermediateXXXwire_922_5,
NOT_intermediateXXXwire_922_6,
NOT_intermediateXXXwire_922_7,
NOT_intermediateXXXwire_795_0,
NOT_intermediateXXXwire_795_1,
NOT_intermediateXXXwire_795_2,
NOT_intermediateXXXwire_795_3,
NOT_intermediateXXXwire_795_4,
NOT_intermediateXXXwire_795_5,
NOT_intermediateXXXwire_795_6,
NOT_intermediateXXXwire_795_7,
NOT_intermediateXXXwire_795_8,
NOT_intermediateXXXwire_795_9,
clk_net_0,
rst_net_0,
start_net_0,
busy_net_0;

pin #(13) pin_0 ({clk, rst, start, func[0], func[1], x[0], x[1], x[2], x[3], x[4], x[5], x[6], x[7]}, {clk_net_0, rst_net_0, start_net_0, func_0, func_1, x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7});

pout #(11) pout_0 ({busy_net_0, resultIPart_0, resultIPart_1, resultFPart_0, resultFPart_1, resultFPart_2, resultFPart_3, resultFPart_4, resultFPart_5, resultFPart_6, resultFPart_7}, {busy, resultIPart[0], resultIPart[1], resultFPart[0], resultFPart[1], resultFPart[2], resultFPart[3], resultFPart[4], resultFPart[5], resultFPart[6], resultFPart[7]});

fanout_n #(2, 0, 0) FANOUT_1 (fourFunc_wire_35, {fourFunc_wire_35_0, fourFunc_wire_35_1});
fanout_n #(2, 0, 0) FANOUT_2 (fourFunc_wire_46, {fourFunc_wire_46_0, fourFunc_wire_46_1});
fanout_n #(3, 0, 0) FANOUT_3 (fourFunc_wire_122, {fourFunc_wire_122_0, fourFunc_wire_122_1, fourFunc_wire_122_2});
fanout_n #(3, 0, 0) FANOUT_4 (fourFunc_wire_133, {fourFunc_wire_133_0, fourFunc_wire_133_1, fourFunc_wire_133_2});
fanout_n #(3, 0, 0) FANOUT_5 (fourFunc_wire_138, {fourFunc_wire_138_0, fourFunc_wire_138_1, fourFunc_wire_138_2});
fanout_n #(3, 0, 0) FANOUT_6 (fourFunc_wire_143, {fourFunc_wire_143_0, fourFunc_wire_143_1, fourFunc_wire_143_2});
fanout_n #(3, 0, 0) FANOUT_7 (fourFunc_wire_148, {fourFunc_wire_148_0, fourFunc_wire_148_1, fourFunc_wire_148_2});
fanout_n #(3, 0, 0) FANOUT_8 (fourFunc_wire_153, {fourFunc_wire_153_0, fourFunc_wire_153_1, fourFunc_wire_153_2});
fanout_n #(3, 0, 0) FANOUT_9 (fourFunc_wire_158, {fourFunc_wire_158_0, fourFunc_wire_158_1, fourFunc_wire_158_2});
fanout_n #(2, 0, 0) FANOUT_10 (fourFunc_wire_184, {fourFunc_wire_184_0, fourFunc_wire_184_1});
fanout_n #(3, 0, 0) FANOUT_11 (fourFunc_wire_166, {fourFunc_wire_166_0, fourFunc_wire_166_1, fourFunc_wire_166_2});
fanout_n #(3, 0, 0) FANOUT_12 (fourFunc_wire_170, {fourFunc_wire_170_0, fourFunc_wire_170_1, fourFunc_wire_170_2});
fanout_n #(3, 0, 0) FANOUT_13 (fourFunc_wire_174, {fourFunc_wire_174_0, fourFunc_wire_174_1, fourFunc_wire_174_2});
fanout_n #(3, 0, 0) FANOUT_14 (fourFunc_wire_178, {fourFunc_wire_178_0, fourFunc_wire_178_1, fourFunc_wire_178_2});
fanout_n #(3, 0, 0) FANOUT_15 (fourFunc_wire_182, {fourFunc_wire_182_0, fourFunc_wire_182_1, fourFunc_wire_182_2});
fanout_n #(3, 0, 0) FANOUT_16 (fourFunc_wire_187, {fourFunc_wire_187_0, fourFunc_wire_187_1, fourFunc_wire_187_2});
fanout_n #(2, 0, 0) FANOUT_17 (fourFunc_wire_213, {fourFunc_wire_213_0, fourFunc_wire_213_1});
fanout_n #(3, 0, 0) FANOUT_18 (fourFunc_wire_195, {fourFunc_wire_195_0, fourFunc_wire_195_1, fourFunc_wire_195_2});
fanout_n #(3, 0, 0) FANOUT_19 (fourFunc_wire_199, {fourFunc_wire_199_0, fourFunc_wire_199_1, fourFunc_wire_199_2});
fanout_n #(3, 0, 0) FANOUT_20 (fourFunc_wire_203, {fourFunc_wire_203_0, fourFunc_wire_203_1, fourFunc_wire_203_2});
fanout_n #(3, 0, 0) FANOUT_21 (fourFunc_wire_207, {fourFunc_wire_207_0, fourFunc_wire_207_1, fourFunc_wire_207_2});
fanout_n #(3, 0, 0) FANOUT_22 (fourFunc_wire_211, {fourFunc_wire_211_0, fourFunc_wire_211_1, fourFunc_wire_211_2});
fanout_n #(3, 0, 0) FANOUT_23 (fourFunc_wire_216, {fourFunc_wire_216_0, fourFunc_wire_216_1, fourFunc_wire_216_2});
fanout_n #(2, 0, 0) FANOUT_24 (fourFunc_wire_242, {fourFunc_wire_242_0, fourFunc_wire_242_1});
fanout_n #(3, 0, 0) FANOUT_25 (fourFunc_wire_224, {fourFunc_wire_224_0, fourFunc_wire_224_1, fourFunc_wire_224_2});
fanout_n #(3, 0, 0) FANOUT_26 (fourFunc_wire_228, {fourFunc_wire_228_0, fourFunc_wire_228_1, fourFunc_wire_228_2});
fanout_n #(3, 0, 0) FANOUT_27 (fourFunc_wire_232, {fourFunc_wire_232_0, fourFunc_wire_232_1, fourFunc_wire_232_2});
fanout_n #(3, 0, 0) FANOUT_28 (fourFunc_wire_236, {fourFunc_wire_236_0, fourFunc_wire_236_1, fourFunc_wire_236_2});
fanout_n #(3, 0, 0) FANOUT_29 (fourFunc_wire_240, {fourFunc_wire_240_0, fourFunc_wire_240_1, fourFunc_wire_240_2});
fanout_n #(3, 0, 0) FANOUT_30 (fourFunc_wire_245, {fourFunc_wire_245_0, fourFunc_wire_245_1, fourFunc_wire_245_2});
fanout_n #(2, 0, 0) FANOUT_31 (fourFunc_wire_271, {fourFunc_wire_271_0, fourFunc_wire_271_1});
fanout_n #(3, 0, 0) FANOUT_32 (fourFunc_wire_253, {fourFunc_wire_253_0, fourFunc_wire_253_1, fourFunc_wire_253_2});
fanout_n #(3, 0, 0) FANOUT_33 (fourFunc_wire_257, {fourFunc_wire_257_0, fourFunc_wire_257_1, fourFunc_wire_257_2});
fanout_n #(3, 0, 0) FANOUT_34 (fourFunc_wire_261, {fourFunc_wire_261_0, fourFunc_wire_261_1, fourFunc_wire_261_2});
fanout_n #(3, 0, 0) FANOUT_35 (fourFunc_wire_265, {fourFunc_wire_265_0, fourFunc_wire_265_1, fourFunc_wire_265_2});
fanout_n #(3, 0, 0) FANOUT_36 (fourFunc_wire_269, {fourFunc_wire_269_0, fourFunc_wire_269_1, fourFunc_wire_269_2});
fanout_n #(3, 0, 0) FANOUT_37 (fourFunc_wire_274, {fourFunc_wire_274_0, fourFunc_wire_274_1, fourFunc_wire_274_2});
fanout_n #(2, 0, 0) FANOUT_38 (fourFunc_wire_299, {fourFunc_wire_299_0, fourFunc_wire_299_1});
fanout_n #(3, 0, 0) FANOUT_39 (fourFunc_wire_285, {fourFunc_wire_285_0, fourFunc_wire_285_1, fourFunc_wire_285_2});
fanout_n #(3, 0, 0) FANOUT_40 (fourFunc_wire_289, {fourFunc_wire_289_0, fourFunc_wire_289_1, fourFunc_wire_289_2});
fanout_n #(3, 0, 0) FANOUT_41 (fourFunc_wire_293, {fourFunc_wire_293_0, fourFunc_wire_293_1, fourFunc_wire_293_2});
fanout_n #(3, 0, 0) FANOUT_42 (fourFunc_wire_297, {fourFunc_wire_297_0, fourFunc_wire_297_1, fourFunc_wire_297_2});
fanout_n #(3, 0, 0) FANOUT_43 (fourFunc_wire_302, {fourFunc_wire_302_0, fourFunc_wire_302_1, fourFunc_wire_302_2});
fanout_n #(2, 0, 0) FANOUT_44 (fourFunc_wire_324, {fourFunc_wire_324_0, fourFunc_wire_324_1});
fanout_n #(2, 0, 0) FANOUT_45 (fourFunc_wire_121, {fourFunc_wire_121_0, fourFunc_wire_121_1});
fanout_n #(2, 0, 0) FANOUT_46 (fourFunc_wire_118, {fourFunc_wire_118_0, fourFunc_wire_118_1});
fanout_n #(2, 0, 0) FANOUT_47 (fourFunc_wire_115, {fourFunc_wire_115_0, fourFunc_wire_115_1});
fanout_n #(2, 0, 0) FANOUT_48 (fourFunc_wire_112, {fourFunc_wire_112_0, fourFunc_wire_112_1});
fanout_n #(2, 0, 0) FANOUT_49 (fourFunc_wire_109, {fourFunc_wire_109_0, fourFunc_wire_109_1});
fanout_n #(2, 0, 0) FANOUT_50 (fourFunc_wire_106, {fourFunc_wire_106_0, fourFunc_wire_106_1});
fanout_n #(2, 0, 0) FANOUT_51 (fourFunc_wire_103, {fourFunc_wire_103_0, fourFunc_wire_103_1});
fanout_n #(2, 0, 0) FANOUT_52 (fourFunc_wire_98, {fourFunc_wire_98_0, fourFunc_wire_98_1});
fanout_n #(2, 0, 0) FANOUT_53 (fourFunc_wire_306, {fourFunc_wire_306_0, fourFunc_wire_306_1});
fanout_n #(2, 0, 0) FANOUT_54 (fourFunc_wire_310, {fourFunc_wire_310_0, fourFunc_wire_310_1});
fanout_n #(2, 0, 0) FANOUT_55 (fourFunc_wire_314, {fourFunc_wire_314_0, fourFunc_wire_314_1});
fanout_n #(2, 0, 0) FANOUT_56 (fourFunc_wire_318, {fourFunc_wire_318_0, fourFunc_wire_318_1});
fanout_n #(2, 0, 0) FANOUT_57 (fourFunc_wire_322, {fourFunc_wire_322_0, fourFunc_wire_322_1});
fanout_n #(2, 0, 0) FANOUT_58 (fourFunc_wire_327, {fourFunc_wire_327_0, fourFunc_wire_327_1});
fanout_n #(3, 0, 0) FANOUT_59 (fourFunc_wire_278, {fourFunc_wire_278_0, fourFunc_wire_278_1, fourFunc_wire_278_2});
fanout_n #(2, 0, 0) FANOUT_60 (fourFunc_wire_124, {fourFunc_wire_124_0, fourFunc_wire_124_1});
fanout_n #(3, 0, 0) FANOUT_61 (fourFunc_wire_307, {fourFunc_wire_307_0, fourFunc_wire_307_1, fourFunc_wire_307_2});
fanout_n #(3, 0, 0) FANOUT_62 (fourFunc_wire_311, {fourFunc_wire_311_0, fourFunc_wire_311_1, fourFunc_wire_311_2});
fanout_n #(3, 0, 0) FANOUT_63 (fourFunc_wire_315, {fourFunc_wire_315_0, fourFunc_wire_315_1, fourFunc_wire_315_2});
fanout_n #(3, 0, 0) FANOUT_64 (fourFunc_wire_319, {fourFunc_wire_319_0, fourFunc_wire_319_1, fourFunc_wire_319_2});
fanout_n #(3, 0, 0) FANOUT_65 (fourFunc_wire_323, {fourFunc_wire_323_0, fourFunc_wire_323_1, fourFunc_wire_323_2});
fanout_n #(2, 0, 0) FANOUT_66 (fourFunc_wire_328, {fourFunc_wire_328_0, fourFunc_wire_328_1});
fanout_n #(2, 0, 0) FANOUT_67 (fourFunc_wire_279, {fourFunc_wire_279_0, fourFunc_wire_279_1});
fanout_n #(2, 0, 0) FANOUT_68 (fourFunc_wire_282, {fourFunc_wire_282_0, fourFunc_wire_282_1});
fanout_n #(2, 0, 0) FANOUT_69 (fourFunc_wire_286, {fourFunc_wire_286_0, fourFunc_wire_286_1});
fanout_n #(2, 0, 0) FANOUT_70 (fourFunc_wire_290, {fourFunc_wire_290_0, fourFunc_wire_290_1});
fanout_n #(2, 0, 0) FANOUT_71 (fourFunc_wire_294, {fourFunc_wire_294_0, fourFunc_wire_294_1});
fanout_n #(2, 0, 0) FANOUT_72 (fourFunc_wire_298, {fourFunc_wire_298_0, fourFunc_wire_298_1});
fanout_n #(2, 0, 0) FANOUT_73 (fourFunc_wire_250, {fourFunc_wire_250_0, fourFunc_wire_250_1});
fanout_n #(2, 0, 0) FANOUT_74 (fourFunc_wire_254, {fourFunc_wire_254_0, fourFunc_wire_254_1});
fanout_n #(2, 0, 0) FANOUT_75 (fourFunc_wire_258, {fourFunc_wire_258_0, fourFunc_wire_258_1});
fanout_n #(2, 0, 0) FANOUT_76 (fourFunc_wire_262, {fourFunc_wire_262_0, fourFunc_wire_262_1});
fanout_n #(2, 0, 0) FANOUT_77 (fourFunc_wire_266, {fourFunc_wire_266_0, fourFunc_wire_266_1});
fanout_n #(2, 0, 0) FANOUT_78 (fourFunc_wire_270, {fourFunc_wire_270_0, fourFunc_wire_270_1});
fanout_n #(2, 0, 0) FANOUT_79 (fourFunc_wire_221, {fourFunc_wire_221_0, fourFunc_wire_221_1});
fanout_n #(2, 0, 0) FANOUT_80 (fourFunc_wire_225, {fourFunc_wire_225_0, fourFunc_wire_225_1});
fanout_n #(2, 0, 0) FANOUT_81 (fourFunc_wire_229, {fourFunc_wire_229_0, fourFunc_wire_229_1});
fanout_n #(2, 0, 0) FANOUT_82 (fourFunc_wire_233, {fourFunc_wire_233_0, fourFunc_wire_233_1});
fanout_n #(2, 0, 0) FANOUT_83 (fourFunc_wire_237, {fourFunc_wire_237_0, fourFunc_wire_237_1});
fanout_n #(2, 0, 0) FANOUT_84 (fourFunc_wire_241, {fourFunc_wire_241_0, fourFunc_wire_241_1});
fanout_n #(2, 0, 0) FANOUT_85 (fourFunc_wire_192, {fourFunc_wire_192_0, fourFunc_wire_192_1});
fanout_n #(2, 0, 0) FANOUT_86 (fourFunc_wire_196, {fourFunc_wire_196_0, fourFunc_wire_196_1});
fanout_n #(2, 0, 0) FANOUT_87 (fourFunc_wire_200, {fourFunc_wire_200_0, fourFunc_wire_200_1});
fanout_n #(2, 0, 0) FANOUT_88 (fourFunc_wire_204, {fourFunc_wire_204_0, fourFunc_wire_204_1});
fanout_n #(2, 0, 0) FANOUT_89 (fourFunc_wire_208, {fourFunc_wire_208_0, fourFunc_wire_208_1});
fanout_n #(2, 0, 0) FANOUT_90 (fourFunc_wire_212, {fourFunc_wire_212_0, fourFunc_wire_212_1});
fanout_n #(2, 0, 0) FANOUT_91 (fourFunc_wire_163, {fourFunc_wire_163_0, fourFunc_wire_163_1});
fanout_n #(2, 0, 0) FANOUT_92 (fourFunc_wire_167, {fourFunc_wire_167_0, fourFunc_wire_167_1});
fanout_n #(2, 0, 0) FANOUT_93 (fourFunc_wire_171, {fourFunc_wire_171_0, fourFunc_wire_171_1});
fanout_n #(2, 0, 0) FANOUT_94 (fourFunc_wire_175, {fourFunc_wire_175_0, fourFunc_wire_175_1});
fanout_n #(2, 0, 0) FANOUT_95 (fourFunc_wire_179, {fourFunc_wire_179_0, fourFunc_wire_179_1});
fanout_n #(2, 0, 0) FANOUT_96 (fourFunc_wire_183, {fourFunc_wire_183_0, fourFunc_wire_183_1});
fanout_n #(2, 0, 0) FANOUT_97 (fourFunc_wire_129, {fourFunc_wire_129_0, fourFunc_wire_129_1});
fanout_n #(2, 0, 0) FANOUT_98 (fourFunc_wire_134, {fourFunc_wire_134_0, fourFunc_wire_134_1});
fanout_n #(2, 0, 0) FANOUT_99 (fourFunc_wire_139, {fourFunc_wire_139_0, fourFunc_wire_139_1});
fanout_n #(2, 0, 0) FANOUT_100 (fourFunc_wire_144, {fourFunc_wire_144_0, fourFunc_wire_144_1});
fanout_n #(2, 0, 0) FANOUT_101 (fourFunc_wire_149, {fourFunc_wire_149_0, fourFunc_wire_149_1});
fanout_n #(2, 0, 0) FANOUT_102 (fourFunc_wire_154, {fourFunc_wire_154_0, fourFunc_wire_154_1});
fanout_n #(3, 0, 0) FANOUT_103 (fourFunc_wire_249, {fourFunc_wire_249_0, fourFunc_wire_249_1, fourFunc_wire_249_2});
fanout_n #(3, 0, 0) FANOUT_104 (fourFunc_wire_220, {fourFunc_wire_220_0, fourFunc_wire_220_1, fourFunc_wire_220_2});
fanout_n #(3, 0, 0) FANOUT_105 (fourFunc_wire_191, {fourFunc_wire_191_0, fourFunc_wire_191_1, fourFunc_wire_191_2});
fanout_n #(3, 0, 0) FANOUT_106 (fourFunc_wire_162, {fourFunc_wire_162_0, fourFunc_wire_162_1, fourFunc_wire_162_2});
fanout_n #(3, 0, 0) FANOUT_107 (fourFunc_wire_128, {fourFunc_wire_128_0, fourFunc_wire_128_1, fourFunc_wire_128_2});
fanout_n #(3, 0, 0) FANOUT_108 (fourFunc_wire_321, {fourFunc_wire_321_0, fourFunc_wire_321_1, fourFunc_wire_321_2});
fanout_n #(3, 0, 0) FANOUT_109 (fourFunc_wire_317, {fourFunc_wire_317_0, fourFunc_wire_317_1, fourFunc_wire_317_2});
fanout_n #(3, 0, 0) FANOUT_110 (fourFunc_wire_313, {fourFunc_wire_313_0, fourFunc_wire_313_1, fourFunc_wire_313_2});
fanout_n #(3, 0, 0) FANOUT_111 (fourFunc_wire_309, {fourFunc_wire_309_0, fourFunc_wire_309_1, fourFunc_wire_309_2});
fanout_n #(3, 0, 0) FANOUT_112 (fourFunc_wire_305, {fourFunc_wire_305_0, fourFunc_wire_305_1, fourFunc_wire_305_2});
fanout_n #(2, 0, 0) FANOUT_113 (fourFunc_wire_123, {fourFunc_wire_123_0, fourFunc_wire_123_1});
fanout_n #(3, 0, 0) FANOUT_114 (fourFunc_wire_296, {fourFunc_wire_296_0, fourFunc_wire_296_1, fourFunc_wire_296_2});
fanout_n #(3, 0, 0) FANOUT_115 (fourFunc_wire_292, {fourFunc_wire_292_0, fourFunc_wire_292_1, fourFunc_wire_292_2});
fanout_n #(3, 0, 0) FANOUT_116 (fourFunc_wire_288, {fourFunc_wire_288_0, fourFunc_wire_288_1, fourFunc_wire_288_2});
fanout_n #(3, 0, 0) FANOUT_117 (fourFunc_wire_284, {fourFunc_wire_284_0, fourFunc_wire_284_1, fourFunc_wire_284_2});
fanout_n #(3, 0, 0) FANOUT_118 (fourFunc_wire_281, {fourFunc_wire_281_0, fourFunc_wire_281_1, fourFunc_wire_281_2});
fanout_n #(3, 0, 0) FANOUT_119 (fourFunc_wire_277, {fourFunc_wire_277_0, fourFunc_wire_277_1, fourFunc_wire_277_2});
fanout_n #(3, 0, 0) FANOUT_120 (fourFunc_wire_268, {fourFunc_wire_268_0, fourFunc_wire_268_1, fourFunc_wire_268_2});
fanout_n #(3, 0, 0) FANOUT_121 (fourFunc_wire_264, {fourFunc_wire_264_0, fourFunc_wire_264_1, fourFunc_wire_264_2});
fanout_n #(3, 0, 0) FANOUT_122 (fourFunc_wire_260, {fourFunc_wire_260_0, fourFunc_wire_260_1, fourFunc_wire_260_2});
fanout_n #(3, 0, 0) FANOUT_123 (fourFunc_wire_256, {fourFunc_wire_256_0, fourFunc_wire_256_1, fourFunc_wire_256_2});
fanout_n #(3, 0, 0) FANOUT_124 (fourFunc_wire_252, {fourFunc_wire_252_0, fourFunc_wire_252_1, fourFunc_wire_252_2});
fanout_n #(3, 0, 0) FANOUT_125 (fourFunc_wire_248, {fourFunc_wire_248_0, fourFunc_wire_248_1, fourFunc_wire_248_2});
fanout_n #(3, 0, 0) FANOUT_126 (fourFunc_wire_239, {fourFunc_wire_239_0, fourFunc_wire_239_1, fourFunc_wire_239_2});
fanout_n #(3, 0, 0) FANOUT_127 (fourFunc_wire_235, {fourFunc_wire_235_0, fourFunc_wire_235_1, fourFunc_wire_235_2});
fanout_n #(3, 0, 0) FANOUT_128 (fourFunc_wire_231, {fourFunc_wire_231_0, fourFunc_wire_231_1, fourFunc_wire_231_2});
fanout_n #(3, 0, 0) FANOUT_129 (fourFunc_wire_227, {fourFunc_wire_227_0, fourFunc_wire_227_1, fourFunc_wire_227_2});
fanout_n #(3, 0, 0) FANOUT_130 (fourFunc_wire_223, {fourFunc_wire_223_0, fourFunc_wire_223_1, fourFunc_wire_223_2});
fanout_n #(3, 0, 0) FANOUT_131 (fourFunc_wire_219, {fourFunc_wire_219_0, fourFunc_wire_219_1, fourFunc_wire_219_2});
fanout_n #(3, 0, 0) FANOUT_132 (fourFunc_wire_210, {fourFunc_wire_210_0, fourFunc_wire_210_1, fourFunc_wire_210_2});
fanout_n #(3, 0, 0) FANOUT_133 (fourFunc_wire_206, {fourFunc_wire_206_0, fourFunc_wire_206_1, fourFunc_wire_206_2});
fanout_n #(3, 0, 0) FANOUT_134 (fourFunc_wire_202, {fourFunc_wire_202_0, fourFunc_wire_202_1, fourFunc_wire_202_2});
fanout_n #(3, 0, 0) FANOUT_135 (fourFunc_wire_198, {fourFunc_wire_198_0, fourFunc_wire_198_1, fourFunc_wire_198_2});
fanout_n #(3, 0, 0) FANOUT_136 (fourFunc_wire_194, {fourFunc_wire_194_0, fourFunc_wire_194_1, fourFunc_wire_194_2});
fanout_n #(3, 0, 0) FANOUT_137 (fourFunc_wire_190, {fourFunc_wire_190_0, fourFunc_wire_190_1, fourFunc_wire_190_2});
fanout_n #(3, 0, 0) FANOUT_138 (fourFunc_wire_181, {fourFunc_wire_181_0, fourFunc_wire_181_1, fourFunc_wire_181_2});
fanout_n #(3, 0, 0) FANOUT_139 (fourFunc_wire_177, {fourFunc_wire_177_0, fourFunc_wire_177_1, fourFunc_wire_177_2});
fanout_n #(3, 0, 0) FANOUT_140 (fourFunc_wire_173, {fourFunc_wire_173_0, fourFunc_wire_173_1, fourFunc_wire_173_2});
fanout_n #(3, 0, 0) FANOUT_141 (fourFunc_wire_169, {fourFunc_wire_169_0, fourFunc_wire_169_1, fourFunc_wire_169_2});
fanout_n #(3, 0, 0) FANOUT_142 (fourFunc_wire_165, {fourFunc_wire_165_0, fourFunc_wire_165_1, fourFunc_wire_165_2});
fanout_n #(3, 0, 0) FANOUT_143 (fourFunc_wire_161, {fourFunc_wire_161_0, fourFunc_wire_161_1, fourFunc_wire_161_2});
fanout_n #(3, 0, 0) FANOUT_144 (fourFunc_wire_152, {fourFunc_wire_152_0, fourFunc_wire_152_1, fourFunc_wire_152_2});
fanout_n #(3, 0, 0) FANOUT_145 (fourFunc_wire_147, {fourFunc_wire_147_0, fourFunc_wire_147_1, fourFunc_wire_147_2});
fanout_n #(3, 0, 0) FANOUT_146 (fourFunc_wire_142, {fourFunc_wire_142_0, fourFunc_wire_142_1, fourFunc_wire_142_2});
fanout_n #(3, 0, 0) FANOUT_147 (fourFunc_wire_137, {fourFunc_wire_137_0, fourFunc_wire_137_1, fourFunc_wire_137_2});
fanout_n #(3, 0, 0) FANOUT_148 (fourFunc_wire_132, {fourFunc_wire_132_0, fourFunc_wire_132_1, fourFunc_wire_132_2});
fanout_n #(3, 0, 0) FANOUT_149 (fourFunc_wire_127, {fourFunc_wire_127_0, fourFunc_wire_127_1, fourFunc_wire_127_2});
fanout_n #(2, 0, 0) FANOUT_150 (fourFunc_wire_93, {fourFunc_wire_93_0, fourFunc_wire_93_1});
fanout_n #(2, 0, 0) FANOUT_151 (fourFunc_wire_88, {fourFunc_wire_88_0, fourFunc_wire_88_1});
fanout_n #(2, 0, 0) FANOUT_152 (fourFunc_wire_83, {fourFunc_wire_83_0, fourFunc_wire_83_1});
fanout_n #(2, 0, 0) FANOUT_153 (fourFunc_wire_78, {fourFunc_wire_78_0, fourFunc_wire_78_1});
fanout_n #(2, 0, 0) FANOUT_154 (fourFunc_wire_73, {fourFunc_wire_73_0, fourFunc_wire_73_1});
fanout_n #(2, 0, 0) FANOUT_155 (fourFunc_wire_68, {fourFunc_wire_68_0, fourFunc_wire_68_1});
fanout_n #(2, 0, 0) FANOUT_156 (fourFunc_wire_63, {fourFunc_wire_63_0, fourFunc_wire_63_1});
fanout_n #(2, 0, 0) FANOUT_157 (fourFunc_wire_60, {fourFunc_wire_60_0, fourFunc_wire_60_1});
fanout_n #(22, 0, 0) FANOUT_158 (fourFunc_wire_551, {fourFunc_wire_551_0, fourFunc_wire_551_1, fourFunc_wire_551_2, fourFunc_wire_551_3, fourFunc_wire_551_4, fourFunc_wire_551_5, fourFunc_wire_551_6, fourFunc_wire_551_7, fourFunc_wire_551_8, fourFunc_wire_551_9, fourFunc_wire_551_10, fourFunc_wire_551_11, fourFunc_wire_551_12, fourFunc_wire_551_13, fourFunc_wire_551_14, fourFunc_wire_551_15, fourFunc_wire_551_16, fourFunc_wire_551_17, fourFunc_wire_551_18, fourFunc_wire_551_19, fourFunc_wire_551_20, fourFunc_wire_551_21});
fanout_n #(11, 0, 0) FANOUT_159 (fourFunc_wire_2, {fourFunc_wire_2_0, fourFunc_wire_2_1, fourFunc_wire_2_2, fourFunc_wire_2_3, fourFunc_wire_2_4, fourFunc_wire_2_5, fourFunc_wire_2_6, fourFunc_wire_2_7, fourFunc_wire_2_8, fourFunc_wire_2_9, fourFunc_wire_2_10});
fanout_n #(11, 0, 0) FANOUT_160 (fourFunc_wire_10, {fourFunc_wire_10_0, fourFunc_wire_10_1, fourFunc_wire_10_2, fourFunc_wire_10_3, fourFunc_wire_10_4, fourFunc_wire_10_5, fourFunc_wire_10_6, fourFunc_wire_10_7, fourFunc_wire_10_8, fourFunc_wire_10_9, fourFunc_wire_10_10});
fanout_n #(9, 0, 0) FANOUT_161 (fourFunc_wire_3, {fourFunc_wire_3_0, fourFunc_wire_3_1, fourFunc_wire_3_2, fourFunc_wire_3_3, fourFunc_wire_3_4, fourFunc_wire_3_5, fourFunc_wire_3_6, fourFunc_wire_3_7, fourFunc_wire_3_8});
fanout_n #(12, 0, 0) FANOUT_162 (fourFunc_wire_8, {fourFunc_wire_8_0, fourFunc_wire_8_1, fourFunc_wire_8_2, fourFunc_wire_8_3, fourFunc_wire_8_4, fourFunc_wire_8_5, fourFunc_wire_8_6, fourFunc_wire_8_7, fourFunc_wire_8_8, fourFunc_wire_8_9, fourFunc_wire_8_10, fourFunc_wire_8_11});
fanout_n #(2, 0, 0) FANOUT_163 (fourFunc_wire_552, {fourFunc_wire_552_0, fourFunc_wire_552_1});
fanout_n #(2, 0, 0) FANOUT_164 (fourFunc_wire_553, {fourFunc_wire_553_0, fourFunc_wire_553_1});
fanout_n #(2, 0, 0) FANOUT_165 (fourFunc_wire_554, {fourFunc_wire_554_0, fourFunc_wire_554_1});
fanout_n #(2, 0, 0) FANOUT_166 (fourFunc_wire_555, {fourFunc_wire_555_0, fourFunc_wire_555_1});
fanout_n #(2, 0, 0) FANOUT_167 (fourFunc_wire_556, {fourFunc_wire_556_0, fourFunc_wire_556_1});
fanout_n #(2, 0, 0) FANOUT_168 (fourFunc_wire_557, {fourFunc_wire_557_0, fourFunc_wire_557_1});
fanout_n #(2, 0, 0) FANOUT_169 (fourFunc_wire_558, {fourFunc_wire_558_0, fourFunc_wire_558_1});
fanout_n #(2, 0, 0) FANOUT_170 (fourFunc_wire_559, {fourFunc_wire_559_0, fourFunc_wire_559_1});
fanout_n #(19, 0, 0) FANOUT_171 (fourFunc_wire_53, {fourFunc_wire_53_0, fourFunc_wire_53_1, fourFunc_wire_53_2, fourFunc_wire_53_3, fourFunc_wire_53_4, fourFunc_wire_53_5, fourFunc_wire_53_6, fourFunc_wire_53_7, fourFunc_wire_53_8, fourFunc_wire_53_9, fourFunc_wire_53_10, fourFunc_wire_53_11, fourFunc_wire_53_12, fourFunc_wire_53_13, fourFunc_wire_53_14, fourFunc_wire_53_15, fourFunc_wire_53_16, fourFunc_wire_53_17, fourFunc_wire_53_18});
fanout_n #(28, 0, 0) FANOUT_172 (fourFunc_wire_95, {fourFunc_wire_95_0, fourFunc_wire_95_1, fourFunc_wire_95_2, fourFunc_wire_95_3, fourFunc_wire_95_4, fourFunc_wire_95_5, fourFunc_wire_95_6, fourFunc_wire_95_7, fourFunc_wire_95_8, fourFunc_wire_95_9, fourFunc_wire_95_10, fourFunc_wire_95_11, fourFunc_wire_95_12, fourFunc_wire_95_13, fourFunc_wire_95_14, fourFunc_wire_95_15, fourFunc_wire_95_16, fourFunc_wire_95_17, fourFunc_wire_95_18, fourFunc_wire_95_19, fourFunc_wire_95_20, fourFunc_wire_95_21, fourFunc_wire_95_22, fourFunc_wire_95_23, fourFunc_wire_95_24, fourFunc_wire_95_25, fourFunc_wire_95_26, fourFunc_wire_95_27});
fanout_n #(15, 0, 0) FANOUT_173 (fourFunc_wire_90, {fourFunc_wire_90_0, fourFunc_wire_90_1, fourFunc_wire_90_2, fourFunc_wire_90_3, fourFunc_wire_90_4, fourFunc_wire_90_5, fourFunc_wire_90_6, fourFunc_wire_90_7, fourFunc_wire_90_8, fourFunc_wire_90_9, fourFunc_wire_90_10, fourFunc_wire_90_11, fourFunc_wire_90_12, fourFunc_wire_90_13, fourFunc_wire_90_14});
fanout_n #(15, 0, 0) FANOUT_174 (fourFunc_wire_85, {fourFunc_wire_85_0, fourFunc_wire_85_1, fourFunc_wire_85_2, fourFunc_wire_85_3, fourFunc_wire_85_4, fourFunc_wire_85_5, fourFunc_wire_85_6, fourFunc_wire_85_7, fourFunc_wire_85_8, fourFunc_wire_85_9, fourFunc_wire_85_10, fourFunc_wire_85_11, fourFunc_wire_85_12, fourFunc_wire_85_13, fourFunc_wire_85_14});
fanout_n #(15, 0, 0) FANOUT_175 (fourFunc_wire_80, {fourFunc_wire_80_0, fourFunc_wire_80_1, fourFunc_wire_80_2, fourFunc_wire_80_3, fourFunc_wire_80_4, fourFunc_wire_80_5, fourFunc_wire_80_6, fourFunc_wire_80_7, fourFunc_wire_80_8, fourFunc_wire_80_9, fourFunc_wire_80_10, fourFunc_wire_80_11, fourFunc_wire_80_12, fourFunc_wire_80_13, fourFunc_wire_80_14});
fanout_n #(15, 0, 0) FANOUT_176 (fourFunc_wire_75, {fourFunc_wire_75_0, fourFunc_wire_75_1, fourFunc_wire_75_2, fourFunc_wire_75_3, fourFunc_wire_75_4, fourFunc_wire_75_5, fourFunc_wire_75_6, fourFunc_wire_75_7, fourFunc_wire_75_8, fourFunc_wire_75_9, fourFunc_wire_75_10, fourFunc_wire_75_11, fourFunc_wire_75_12, fourFunc_wire_75_13, fourFunc_wire_75_14});
fanout_n #(15, 0, 0) FANOUT_177 (fourFunc_wire_70, {fourFunc_wire_70_0, fourFunc_wire_70_1, fourFunc_wire_70_2, fourFunc_wire_70_3, fourFunc_wire_70_4, fourFunc_wire_70_5, fourFunc_wire_70_6, fourFunc_wire_70_7, fourFunc_wire_70_8, fourFunc_wire_70_9, fourFunc_wire_70_10, fourFunc_wire_70_11, fourFunc_wire_70_12, fourFunc_wire_70_13, fourFunc_wire_70_14});
fanout_n #(15, 0, 0) FANOUT_178 (fourFunc_wire_65, {fourFunc_wire_65_0, fourFunc_wire_65_1, fourFunc_wire_65_2, fourFunc_wire_65_3, fourFunc_wire_65_4, fourFunc_wire_65_5, fourFunc_wire_65_6, fourFunc_wire_65_7, fourFunc_wire_65_8, fourFunc_wire_65_9, fourFunc_wire_65_10, fourFunc_wire_65_11, fourFunc_wire_65_12, fourFunc_wire_65_13, fourFunc_wire_65_14});
fanout_n #(6, 0, 0) FANOUT_179 (fourFunc_wire_54, {fourFunc_wire_54_0, fourFunc_wire_54_1, fourFunc_wire_54_2, fourFunc_wire_54_3, fourFunc_wire_54_4, fourFunc_wire_54_5});
fanout_n #(8, 0, 0) FANOUT_180 (fourFunc_wire_94, {fourFunc_wire_94_0, fourFunc_wire_94_1, fourFunc_wire_94_2, fourFunc_wire_94_3, fourFunc_wire_94_4, fourFunc_wire_94_5, fourFunc_wire_94_6, fourFunc_wire_94_7});
fanout_n #(8, 0, 0) FANOUT_181 (fourFunc_wire_89, {fourFunc_wire_89_0, fourFunc_wire_89_1, fourFunc_wire_89_2, fourFunc_wire_89_3, fourFunc_wire_89_4, fourFunc_wire_89_5, fourFunc_wire_89_6, fourFunc_wire_89_7});
fanout_n #(8, 0, 0) FANOUT_182 (fourFunc_wire_84, {fourFunc_wire_84_0, fourFunc_wire_84_1, fourFunc_wire_84_2, fourFunc_wire_84_3, fourFunc_wire_84_4, fourFunc_wire_84_5, fourFunc_wire_84_6, fourFunc_wire_84_7});
fanout_n #(8, 0, 0) FANOUT_183 (fourFunc_wire_79, {fourFunc_wire_79_0, fourFunc_wire_79_1, fourFunc_wire_79_2, fourFunc_wire_79_3, fourFunc_wire_79_4, fourFunc_wire_79_5, fourFunc_wire_79_6, fourFunc_wire_79_7});
fanout_n #(8, 0, 0) FANOUT_184 (fourFunc_wire_74, {fourFunc_wire_74_0, fourFunc_wire_74_1, fourFunc_wire_74_2, fourFunc_wire_74_3, fourFunc_wire_74_4, fourFunc_wire_74_5, fourFunc_wire_74_6, fourFunc_wire_74_7});
fanout_n #(8, 0, 0) FANOUT_185 (fourFunc_wire_69, {fourFunc_wire_69_0, fourFunc_wire_69_1, fourFunc_wire_69_2, fourFunc_wire_69_3, fourFunc_wire_69_4, fourFunc_wire_69_5, fourFunc_wire_69_6, fourFunc_wire_69_7});
fanout_n #(8, 0, 0) FANOUT_186 (fourFunc_wire_64, {fourFunc_wire_64_0, fourFunc_wire_64_1, fourFunc_wire_64_2, fourFunc_wire_64_3, fourFunc_wire_64_4, fourFunc_wire_64_5, fourFunc_wire_64_6, fourFunc_wire_64_7});
fanout_n #(6, 0, 0) FANOUT_187 (fourFunc_wire_59, {fourFunc_wire_59_0, fourFunc_wire_59_1, fourFunc_wire_59_2, fourFunc_wire_59_3, fourFunc_wire_59_4, fourFunc_wire_59_5});
fanout_n #(4, 0, 0) FANOUT_188 (fourFunc_wire_56, {fourFunc_wire_56_0, fourFunc_wire_56_1, fourFunc_wire_56_2, fourFunc_wire_56_3});
fanout_n #(2, 0, 0) FANOUT_189 (fourFunc_wire_582, {fourFunc_wire_582_0, fourFunc_wire_582_1});
fanout_n #(4, 0, 0) FANOUT_190 (fourFunc_wire_588, {fourFunc_wire_588_0, fourFunc_wire_588_1, fourFunc_wire_588_2, fourFunc_wire_588_3});
fanout_n #(5, 0, 0) FANOUT_191 (fourFunc_wire_589, {fourFunc_wire_589_0, fourFunc_wire_589_1, fourFunc_wire_589_2, fourFunc_wire_589_3, fourFunc_wire_589_4});
fanout_n #(3, 0, 0) FANOUT_192 (fourFunc_wire_590, {fourFunc_wire_590_0, fourFunc_wire_590_1, fourFunc_wire_590_2});
fanout_n #(18, 0, 0) FANOUT_193 (fourFunc_wire_586, {fourFunc_wire_586_0, fourFunc_wire_586_1, fourFunc_wire_586_2, fourFunc_wire_586_3, fourFunc_wire_586_4, fourFunc_wire_586_5, fourFunc_wire_586_6, fourFunc_wire_586_7, fourFunc_wire_586_8, fourFunc_wire_586_9, fourFunc_wire_586_10, fourFunc_wire_586_11, fourFunc_wire_586_12, fourFunc_wire_586_13, fourFunc_wire_586_14, fourFunc_wire_586_15, fourFunc_wire_586_16, fourFunc_wire_586_17});
fanout_n #(5, 0, 0) FANOUT_194 (fourFunc_wire_581, {fourFunc_wire_581_0, fourFunc_wire_581_1, fourFunc_wire_581_2, fourFunc_wire_581_3, fourFunc_wire_581_4});
fanout_n #(32, 0, 0) FANOUT_195 (fourFunc_wire_599, {fourFunc_wire_599_0, fourFunc_wire_599_1, fourFunc_wire_599_2, fourFunc_wire_599_3, fourFunc_wire_599_4, fourFunc_wire_599_5, fourFunc_wire_599_6, fourFunc_wire_599_7, fourFunc_wire_599_8, fourFunc_wire_599_9, fourFunc_wire_599_10, fourFunc_wire_599_11, fourFunc_wire_599_12, fourFunc_wire_599_13, fourFunc_wire_599_14, fourFunc_wire_599_15, fourFunc_wire_599_16, fourFunc_wire_599_17, fourFunc_wire_599_18, fourFunc_wire_599_19, fourFunc_wire_599_20, fourFunc_wire_599_21, fourFunc_wire_599_22, fourFunc_wire_599_23, fourFunc_wire_599_24, fourFunc_wire_599_25, fourFunc_wire_599_26, fourFunc_wire_599_27, fourFunc_wire_599_28, fourFunc_wire_599_29, fourFunc_wire_599_30, fourFunc_wire_599_31});
fanout_n #(2, 0, 0) FANOUT_196 (fourFunc_wire_50, {fourFunc_wire_50_0, fourFunc_wire_50_1});
fanout_n #(2, 0, 0) FANOUT_197 (fourFunc_wire_605, {fourFunc_wire_605_0, fourFunc_wire_605_1});
fanout_n #(4, 0, 0) FANOUT_198 (fourFunc_wire_609, {fourFunc_wire_609_0, fourFunc_wire_609_1, fourFunc_wire_609_2, fourFunc_wire_609_3});
fanout_n #(13, 0, 0) FANOUT_199 (fourFunc_wire_608, {fourFunc_wire_608_0, fourFunc_wire_608_1, fourFunc_wire_608_2, fourFunc_wire_608_3, fourFunc_wire_608_4, fourFunc_wire_608_5, fourFunc_wire_608_6, fourFunc_wire_608_7, fourFunc_wire_608_8, fourFunc_wire_608_9, fourFunc_wire_608_10, fourFunc_wire_608_11, fourFunc_wire_608_12});
fanout_n #(40, 0, 0) FANOUT_200 (fourFunc_wire_604, {fourFunc_wire_604_0, fourFunc_wire_604_1, fourFunc_wire_604_2, fourFunc_wire_604_3, fourFunc_wire_604_4, fourFunc_wire_604_5, fourFunc_wire_604_6, fourFunc_wire_604_7, fourFunc_wire_604_8, fourFunc_wire_604_9, fourFunc_wire_604_10, fourFunc_wire_604_11, fourFunc_wire_604_12, fourFunc_wire_604_13, fourFunc_wire_604_14, fourFunc_wire_604_15, fourFunc_wire_604_16, fourFunc_wire_604_17, fourFunc_wire_604_18, fourFunc_wire_604_19, fourFunc_wire_604_20, fourFunc_wire_604_21, fourFunc_wire_604_22, fourFunc_wire_604_23, fourFunc_wire_604_24, fourFunc_wire_604_25, fourFunc_wire_604_26, fourFunc_wire_604_27, fourFunc_wire_604_28, fourFunc_wire_604_29, fourFunc_wire_604_30, fourFunc_wire_604_31, fourFunc_wire_604_32, fourFunc_wire_604_33, fourFunc_wire_604_34, fourFunc_wire_604_35, fourFunc_wire_604_36, fourFunc_wire_604_37, fourFunc_wire_604_38, fourFunc_wire_604_39});
fanout_n #(11, 0, 0) FANOUT_201 (fourFunc_wire_648, {fourFunc_wire_648_0, fourFunc_wire_648_1, fourFunc_wire_648_2, fourFunc_wire_648_3, fourFunc_wire_648_4, fourFunc_wire_648_5, fourFunc_wire_648_6, fourFunc_wire_648_7, fourFunc_wire_648_8, fourFunc_wire_648_9, fourFunc_wire_648_10});
fanout_n #(8, 0, 0) FANOUT_202 (fourFunc_wire_434, {fourFunc_wire_434_0, fourFunc_wire_434_1, fourFunc_wire_434_2, fourFunc_wire_434_3, fourFunc_wire_434_4, fourFunc_wire_434_5, fourFunc_wire_434_6, fourFunc_wire_434_7});
fanout_n #(9, 0, 0) FANOUT_203 (fourFunc_wire_446, {fourFunc_wire_446_0, fourFunc_wire_446_1, fourFunc_wire_446_2, fourFunc_wire_446_3, fourFunc_wire_446_4, fourFunc_wire_446_5, fourFunc_wire_446_6, fourFunc_wire_446_7, fourFunc_wire_446_8});
fanout_n #(9, 0, 0) FANOUT_204 (fourFunc_wire_350, {fourFunc_wire_350_0, fourFunc_wire_350_1, fourFunc_wire_350_2, fourFunc_wire_350_3, fourFunc_wire_350_4, fourFunc_wire_350_5, fourFunc_wire_350_6, fourFunc_wire_350_7, fourFunc_wire_350_8});
fanout_n #(9, 0, 0) FANOUT_205 (fourFunc_wire_364, {fourFunc_wire_364_0, fourFunc_wire_364_1, fourFunc_wire_364_2, fourFunc_wire_364_3, fourFunc_wire_364_4, fourFunc_wire_364_5, fourFunc_wire_364_6, fourFunc_wire_364_7, fourFunc_wire_364_8});
fanout_n #(9, 0, 0) FANOUT_206 (fourFunc_wire_378, {fourFunc_wire_378_0, fourFunc_wire_378_1, fourFunc_wire_378_2, fourFunc_wire_378_3, fourFunc_wire_378_4, fourFunc_wire_378_5, fourFunc_wire_378_6, fourFunc_wire_378_7, fourFunc_wire_378_8});
fanout_n #(9, 0, 0) FANOUT_207 (fourFunc_wire_392, {fourFunc_wire_392_0, fourFunc_wire_392_1, fourFunc_wire_392_2, fourFunc_wire_392_3, fourFunc_wire_392_4, fourFunc_wire_392_5, fourFunc_wire_392_6, fourFunc_wire_392_7, fourFunc_wire_392_8});
fanout_n #(9, 0, 0) FANOUT_208 (fourFunc_wire_406, {fourFunc_wire_406_0, fourFunc_wire_406_1, fourFunc_wire_406_2, fourFunc_wire_406_3, fourFunc_wire_406_4, fourFunc_wire_406_5, fourFunc_wire_406_6, fourFunc_wire_406_7, fourFunc_wire_406_8});
fanout_n #(9, 0, 0) FANOUT_209 (fourFunc_wire_420, {fourFunc_wire_420_0, fourFunc_wire_420_1, fourFunc_wire_420_2, fourFunc_wire_420_3, fourFunc_wire_420_4, fourFunc_wire_420_5, fourFunc_wire_420_6, fourFunc_wire_420_7, fourFunc_wire_420_8});
fanout_n #(9, 0, 0) FANOUT_210 (fourFunc_wire_717, {fourFunc_wire_717_0, fourFunc_wire_717_1, fourFunc_wire_717_2, fourFunc_wire_717_3, fourFunc_wire_717_4, fourFunc_wire_717_5, fourFunc_wire_717_6, fourFunc_wire_717_7, fourFunc_wire_717_8});
fanout_n #(24, 0, 0) FANOUT_211 (fourFunc_wire_9, {fourFunc_wire_9_0, fourFunc_wire_9_1, fourFunc_wire_9_2, fourFunc_wire_9_3, fourFunc_wire_9_4, fourFunc_wire_9_5, fourFunc_wire_9_6, fourFunc_wire_9_7, fourFunc_wire_9_8, fourFunc_wire_9_9, fourFunc_wire_9_10, fourFunc_wire_9_11, fourFunc_wire_9_12, fourFunc_wire_9_13, fourFunc_wire_9_14, fourFunc_wire_9_15, fourFunc_wire_9_16, fourFunc_wire_9_17, fourFunc_wire_9_18, fourFunc_wire_9_19, fourFunc_wire_9_20, fourFunc_wire_9_21, fourFunc_wire_9_22, fourFunc_wire_9_23});
fanout_n #(6, 0, 0) FANOUT_212 (fourFunc_wire_598, {fourFunc_wire_598_0, fourFunc_wire_598_1, fourFunc_wire_598_2, fourFunc_wire_598_3, fourFunc_wire_598_4, fourFunc_wire_598_5});
fanout_n #(3, 0, 0) FANOUT_213 (fourFunc_wire_641, {fourFunc_wire_641_0, fourFunc_wire_641_1, fourFunc_wire_641_2});
fanout_n #(3, 0, 0) FANOUT_214 (fourFunc_wire_626, {fourFunc_wire_626_0, fourFunc_wire_626_1, fourFunc_wire_626_2});
fanout_n #(3, 0, 0) FANOUT_215 (fourFunc_wire_628, {fourFunc_wire_628_0, fourFunc_wire_628_1, fourFunc_wire_628_2});
fanout_n #(3, 0, 0) FANOUT_216 (fourFunc_wire_630, {fourFunc_wire_630_0, fourFunc_wire_630_1, fourFunc_wire_630_2});
fanout_n #(3, 0, 0) FANOUT_217 (fourFunc_wire_634, {fourFunc_wire_634_0, fourFunc_wire_634_1, fourFunc_wire_634_2});
fanout_n #(3, 0, 0) FANOUT_218 (fourFunc_wire_636, {fourFunc_wire_636_0, fourFunc_wire_636_1, fourFunc_wire_636_2});
fanout_n #(3, 0, 0) FANOUT_219 (fourFunc_wire_632, {fourFunc_wire_632_0, fourFunc_wire_632_1, fourFunc_wire_632_2});
fanout_n #(3, 0, 0) FANOUT_220 (fourFunc_wire_638, {fourFunc_wire_638_0, fourFunc_wire_638_1, fourFunc_wire_638_2});
fanout_n #(3, 0, 0) FANOUT_221 (fourFunc_wire_640, {fourFunc_wire_640_0, fourFunc_wire_640_1, fourFunc_wire_640_2});
fanout_n #(3, 0, 0) FANOUT_222 (NOT_intermediateXXXwire_690, {NOT_intermediateXXXwire_690_0, NOT_intermediateXXXwire_690_1, NOT_intermediateXXXwire_690_2});
fanout_n #(8, 0, 0) FANOUT_223 (NOT_intermediateXXXwire_697, {NOT_intermediateXXXwire_697_0, NOT_intermediateXXXwire_697_1, NOT_intermediateXXXwire_697_2, NOT_intermediateXXXwire_697_3, NOT_intermediateXXXwire_697_4, NOT_intermediateXXXwire_697_5, NOT_intermediateXXXwire_697_6, NOT_intermediateXXXwire_697_7});
fanout_n #(8, 0, 0) FANOUT_224 (NOT_intermediateXXXwire_922, {NOT_intermediateXXXwire_922_0, NOT_intermediateXXXwire_922_1, NOT_intermediateXXXwire_922_2, NOT_intermediateXXXwire_922_3, NOT_intermediateXXXwire_922_4, NOT_intermediateXXXwire_922_5, NOT_intermediateXXXwire_922_6, NOT_intermediateXXXwire_922_7});
fanout_n #(10, 0, 0) FANOUT_225 (NOT_intermediateXXXwire_795, {NOT_intermediateXXXwire_795_0, NOT_intermediateXXXwire_795_1, NOT_intermediateXXXwire_795_2, NOT_intermediateXXXwire_795_3, NOT_intermediateXXXwire_795_4, NOT_intermediateXXXwire_795_5, NOT_intermediateXXXwire_795_6, NOT_intermediateXXXwire_795_7, NOT_intermediateXXXwire_795_8, NOT_intermediateXXXwire_795_9});


and_n #(2, 0, 0) AND_1 (fourFunc_wire_1, {fourFunc_wire_2_0, fourFunc_wire_3_0});
and_n #(3, 0, 0) AND_2 (fourFunc_wire_4, {fourFunc_wire_1, fourFunc_wire_5, fourFunc_wire_6});
notg #(0, 0) NOT_1 (fourFunc_wire_7, fourFunc_wire_8_0);
and_n #(2, 0, 0) AND_3 (fourFunc_wire_6, {fourFunc_wire_7, fourFunc_wire_9_0});
notg #(0, 0) NOT_2 (fourFunc_wire_5, fourFunc_wire_10_0);
and_n #(2, 0, 0) AND_4 (fourFunc_wire_11, {fourFunc_wire_2_1, fourFunc_wire_8_1});
and_n #(3, 0, 0) AND_5 (fourFunc_wire_12, {fourFunc_wire_11, fourFunc_wire_13, fourFunc_wire_14});
notg #(0, 0) NOT_3 (fourFunc_wire_15, fourFunc_wire_3_1);
and_n #(2, 0, 0) AND_6 (fourFunc_wire_14, {fourFunc_wire_15, fourFunc_wire_9_1});
notg #(0, 0) NOT_4 (fourFunc_wire_13, fourFunc_wire_10_1);
and_n #(2, 0, 0) AND_7 (fourFunc_wire_16, {fourFunc_wire_2_2, fourFunc_wire_9_2});
and_n #(3, 0, 0) AND_8 (fourFunc_wire_17, {fourFunc_wire_16, fourFunc_wire_18, fourFunc_wire_19});
nor_n #(2, 0, 0) NOR_1 (fourFunc_wire_19, {fourFunc_wire_8_2, fourFunc_wire_3_2});
notg #(0, 0) NOT_5 (fourFunc_wire_18, fourFunc_wire_10_2);
notg #(0, 0) NOT_6 (fourFunc_wire_20, fourFunc_wire_2_3);
notg #(0, 0) NOT_7 (fourFunc_wire_21, fourFunc_wire_2_4);
notg #(0, 0) NOT_8 (fourFunc_wire_22, fourFunc_wire_2_5);
or_n #(2, 0, 0) OR_1 (fourFunc_wire_23, {fourFunc_wire_2_6, fourFunc_wire_24});
and_n #(3, 0, 0) AND_9 (fourFunc_wire_25, {fourFunc_wire_8_3, fourFunc_wire_20, fourFunc_wire_26});
or_n #(2, 0, 0) OR_2 (fourFunc_wire_27, {fourFunc_wire_8_4, fourFunc_wire_28});
and_n #(2, 0, 0) AND_10 (fourFunc_wire_29, {fourFunc_wire_8_5, fourFunc_wire_30});
or_n #(2, 0, 0) OR_3 (fourFunc_wire_31, {fourFunc_wire_8_6, fourFunc_wire_32});
or_n #(2, 0, 0) OR_4 (fourFunc_wire_33, {fourFunc_wire_3_3, fourFunc_wire_10_3});
notg #(0, 0) NOT_9 (fourFunc_wire_34, fourFunc_wire_3_4);
or_n #(3, 0, 0) OR_5 (fourFunc_wire_35, {fourFunc_wire_10_4, fourFunc_wire_34, fourFunc_wire_36});
or_n #(2, 0, 0) OR_6 (fourFunc_wire_37, {fourFunc_wire_10_5, fourFunc_wire_38});
notg #(0, 0) NOT_10 (fourFunc_wire_39, fourFunc_wire_9_3);
notg #(0, 0) NOT_11 (fourFunc_wire_36, fourFunc_wire_9_4);
notg #(0, 0) NOT_12 (fourFunc_wire_38, fourFunc_wire_9_5);
and_n #(2, 0, 0) AND_11 (fourFunc_wire_40, {fourFunc_wire_41, fourFunc_wire_23});
and_n #(3, 0, 0) AND_12 (fourFunc_wire_42, {fourFunc_wire_21, fourFunc_wire_27, fourFunc_wire_43});
or_n #(2, 0, 0) OR_7 (fourFunc_wire_41, {fourFunc_wire_29, fourFunc_wire_22});
nor_n #(2, 0, 0) NOR_2 (fourFunc_wire_32, {fourFunc_wire_44, fourFunc_wire_3_5});
nand_n #(2, 0, 0) NAND_1 (fourFunc_wire_45, {fourFunc_wire_37, fourFunc_wire_8_7});
and_n #(2, 0, 0) AND_13 (fourFunc_wire_24, {fourFunc_wire_45, fourFunc_wire_31});
nand_n #(2, 0, 0) NAND_2 (fourFunc_wire_44, {fourFunc_wire_10_6, fourFunc_wire_9_6});
notg #(0, 0) NOT_13 (fourFunc_wire_30, fourFunc_wire_35_0);
notg #(0, 0) NOT_14 (fourFunc_wire_28, fourFunc_wire_35_1);
or_n #(2, 0, 0) OR_8 (fourFunc_wire_46, {fourFunc_wire_33, fourFunc_wire_39});
nand_n #(2, 0, 0) NAND_3 (fourFunc_wire_43, {fourFunc_wire_8_8, fourFunc_wire_46_0});
notg #(0, 0) NOT_15 (fourFunc_wire_26, fourFunc_wire_46_1);
xor_n #(2, 0, 0) XOR_1 (fourFunc_wire_47, {fourFunc_wire_48, fourFunc_wire_10_7});
xor_n #(2, 0, 0) XOR_2 (fourFunc_wire_49, {fourFunc_wire_50_0, fourFunc_wire_3_6});
xor_n #(2, 0, 0) XOR_3 (fourFunc_wire_51, {fourFunc_wire_2_7, fourFunc_wire_8_9});
xnor_n #(2, 0, 0) XNOR_1 (fourFunc_wire_52, {fourFunc_wire_53_0, fourFunc_wire_54_0});
xnor_n #(2, 0, 0) XNOR_2 (fourFunc_wire_55, {fourFunc_wire_56_0, fourFunc_wire_57});
xnor_n #(2, 0, 0) XNOR_3 (fourFunc_wire_58, {fourFunc_wire_59_0, fourFunc_wire_60_0});
xor_n #(2, 0, 0) XOR_4 (fourFunc_wire_61, {fourFunc_wire_62, fourFunc_wire_63_0});
xnor_n #(2, 0, 0) XNOR_4 (fourFunc_wire_62, {fourFunc_wire_64_0, fourFunc_wire_65_0});
xor_n #(2, 0, 0) XOR_5 (fourFunc_wire_66, {fourFunc_wire_67, fourFunc_wire_68_0});
xnor_n #(2, 0, 0) XNOR_5 (fourFunc_wire_67, {fourFunc_wire_69_0, fourFunc_wire_70_0});
xor_n #(2, 0, 0) XOR_6 (fourFunc_wire_71, {fourFunc_wire_72, fourFunc_wire_73_0});
xnor_n #(2, 0, 0) XNOR_6 (fourFunc_wire_72, {fourFunc_wire_74_0, fourFunc_wire_75_0});
xor_n #(2, 0, 0) XOR_7 (fourFunc_wire_76, {fourFunc_wire_77, fourFunc_wire_78_0});
xnor_n #(2, 0, 0) XNOR_7 (fourFunc_wire_77, {fourFunc_wire_79_0, fourFunc_wire_80_0});
xor_n #(2, 0, 0) XOR_8 (fourFunc_wire_81, {fourFunc_wire_82, fourFunc_wire_83_0});
xnor_n #(2, 0, 0) XNOR_8 (fourFunc_wire_82, {fourFunc_wire_84_0, fourFunc_wire_85_0});
xor_n #(2, 0, 0) XOR_9 (fourFunc_wire_86, {fourFunc_wire_87, fourFunc_wire_88_0});
xnor_n #(2, 0, 0) XNOR_9 (fourFunc_wire_87, {fourFunc_wire_89_0, fourFunc_wire_90_0});
xor_n #(2, 0, 0) XOR_10 (fourFunc_wire_91, {fourFunc_wire_92, fourFunc_wire_93_0});
xnor_n #(2, 0, 0) XNOR_10 (fourFunc_wire_92, {fourFunc_wire_94_0, fourFunc_wire_95_0});
xor_n #(2, 0, 0) XOR_11 (fourFunc_wire_96, {fourFunc_wire_54_1, fourFunc_wire_53_1});
xor_n #(2, 0, 0) XOR_12 (fourFunc_wire_97, {fourFunc_wire_98_0, fourFunc_wire_59_1});
xor_n #(2, 0, 0) XOR_13 (fourFunc_wire_99, {fourFunc_wire_100, fourFunc_wire_56_1});
xor_n #(2, 0, 0) XOR_14 (fourFunc_wire_101, {fourFunc_wire_102, fourFunc_wire_103_0});
xor_n #(2, 0, 0) XOR_15 (fourFunc_wire_102, {fourFunc_wire_65_1, fourFunc_wire_64_1});
xor_n #(2, 0, 0) XOR_16 (fourFunc_wire_104, {fourFunc_wire_105, fourFunc_wire_106_0});
xor_n #(2, 0, 0) XOR_17 (fourFunc_wire_105, {fourFunc_wire_70_1, fourFunc_wire_69_1});
xor_n #(2, 0, 0) XOR_18 (fourFunc_wire_107, {fourFunc_wire_108, fourFunc_wire_109_0});
xor_n #(2, 0, 0) XOR_19 (fourFunc_wire_108, {fourFunc_wire_75_1, fourFunc_wire_74_1});
xor_n #(2, 0, 0) XOR_20 (fourFunc_wire_110, {fourFunc_wire_111, fourFunc_wire_112_0});
xor_n #(2, 0, 0) XOR_21 (fourFunc_wire_111, {fourFunc_wire_80_1, fourFunc_wire_79_1});
xor_n #(2, 0, 0) XOR_22 (fourFunc_wire_113, {fourFunc_wire_114, fourFunc_wire_115_0});
xor_n #(2, 0, 0) XOR_23 (fourFunc_wire_114, {fourFunc_wire_85_1, fourFunc_wire_84_1});
xor_n #(2, 0, 0) XOR_24 (fourFunc_wire_116, {fourFunc_wire_117, fourFunc_wire_118_0});
xor_n #(2, 0, 0) XOR_25 (fourFunc_wire_117, {fourFunc_wire_90_1, fourFunc_wire_89_1});
xor_n #(2, 0, 0) XOR_26 (fourFunc_wire_119, {fourFunc_wire_120, fourFunc_wire_121_0});
xor_n #(2, 0, 0) XOR_27 (fourFunc_wire_120, {fourFunc_wire_95_1, fourFunc_wire_94_1});
xor_n #(2, 0, 0) XOR_28 (fourFunc_wire_122, {fourFunc_wire_123_0, fourFunc_wire_124_0});
xor_n #(2, 0, 0) XOR_29 (fourFunc_wire_125, {fourFunc_wire_126, fourFunc_wire_127_0});
xor_n #(2, 0, 0) XOR_30 (fourFunc_wire_126, {fourFunc_wire_128_0, fourFunc_wire_129_0});
xor_n #(2, 0, 0) XOR_31 (fourFunc_wire_130, {fourFunc_wire_131, fourFunc_wire_132_0});
xor_n #(2, 0, 0) XOR_32 (fourFunc_wire_131, {fourFunc_wire_133_0, fourFunc_wire_134_0});
xor_n #(2, 0, 0) XOR_33 (fourFunc_wire_135, {fourFunc_wire_136, fourFunc_wire_137_0});
xor_n #(2, 0, 0) XOR_34 (fourFunc_wire_136, {fourFunc_wire_138_0, fourFunc_wire_139_0});
xor_n #(2, 0, 0) XOR_35 (fourFunc_wire_140, {fourFunc_wire_141, fourFunc_wire_142_0});
xor_n #(2, 0, 0) XOR_36 (fourFunc_wire_141, {fourFunc_wire_143_0, fourFunc_wire_144_0});
xor_n #(2, 0, 0) XOR_37 (fourFunc_wire_145, {fourFunc_wire_146, fourFunc_wire_147_0});
xor_n #(2, 0, 0) XOR_38 (fourFunc_wire_146, {fourFunc_wire_148_0, fourFunc_wire_149_0});
xor_n #(2, 0, 0) XOR_39 (fourFunc_wire_150, {fourFunc_wire_151, fourFunc_wire_152_0});
xor_n #(2, 0, 0) XOR_40 (fourFunc_wire_151, {fourFunc_wire_153_0, fourFunc_wire_154_0});
xor_n #(2, 0, 0) XOR_41 (fourFunc_wire_155, {fourFunc_wire_156, fourFunc_wire_157});
xor_n #(2, 0, 0) XOR_42 (fourFunc_wire_156, {fourFunc_wire_158_0, fourFunc_wire_159});
xor_n #(2, 0, 0) XOR_43 (fourFunc_wire_133, {fourFunc_wire_160, fourFunc_wire_161_0});
xor_n #(2, 0, 0) XOR_44 (fourFunc_wire_160, {fourFunc_wire_162_0, fourFunc_wire_163_0});
xor_n #(2, 0, 0) XOR_45 (fourFunc_wire_138, {fourFunc_wire_164, fourFunc_wire_165_0});
xor_n #(2, 0, 0) XOR_46 (fourFunc_wire_164, {fourFunc_wire_166_0, fourFunc_wire_167_0});
xor_n #(2, 0, 0) XOR_47 (fourFunc_wire_143, {fourFunc_wire_168, fourFunc_wire_169_0});
xor_n #(2, 0, 0) XOR_48 (fourFunc_wire_168, {fourFunc_wire_170_0, fourFunc_wire_171_0});
xor_n #(2, 0, 0) XOR_49 (fourFunc_wire_148, {fourFunc_wire_172, fourFunc_wire_173_0});
xor_n #(2, 0, 0) XOR_50 (fourFunc_wire_172, {fourFunc_wire_174_0, fourFunc_wire_175_0});
xor_n #(2, 0, 0) XOR_51 (fourFunc_wire_153, {fourFunc_wire_176, fourFunc_wire_177_0});
xor_n #(2, 0, 0) XOR_52 (fourFunc_wire_176, {fourFunc_wire_178_0, fourFunc_wire_179_0});
xor_n #(2, 0, 0) XOR_53 (fourFunc_wire_158, {fourFunc_wire_180, fourFunc_wire_181_0});
xor_n #(2, 0, 0) XOR_54 (fourFunc_wire_180, {fourFunc_wire_182_0, fourFunc_wire_183_0});
xor_n #(2, 0, 0) XOR_55 (fourFunc_wire_184, {fourFunc_wire_185, fourFunc_wire_186});
xor_n #(2, 0, 0) XOR_56 (fourFunc_wire_185, {fourFunc_wire_187_0, fourFunc_wire_188});
xor_n #(2, 0, 0) XOR_57 (fourFunc_wire_166, {fourFunc_wire_189, fourFunc_wire_190_0});
xor_n #(2, 0, 0) XOR_58 (fourFunc_wire_189, {fourFunc_wire_191_0, fourFunc_wire_192_0});
xor_n #(2, 0, 0) XOR_59 (fourFunc_wire_170, {fourFunc_wire_193, fourFunc_wire_194_0});
xor_n #(2, 0, 0) XOR_60 (fourFunc_wire_193, {fourFunc_wire_195_0, fourFunc_wire_196_0});
xor_n #(2, 0, 0) XOR_61 (fourFunc_wire_174, {fourFunc_wire_197, fourFunc_wire_198_0});
xor_n #(2, 0, 0) XOR_62 (fourFunc_wire_197, {fourFunc_wire_199_0, fourFunc_wire_200_0});
xor_n #(2, 0, 0) XOR_63 (fourFunc_wire_178, {fourFunc_wire_201, fourFunc_wire_202_0});
xor_n #(2, 0, 0) XOR_64 (fourFunc_wire_201, {fourFunc_wire_203_0, fourFunc_wire_204_0});
xor_n #(2, 0, 0) XOR_65 (fourFunc_wire_182, {fourFunc_wire_205, fourFunc_wire_206_0});
xor_n #(2, 0, 0) XOR_66 (fourFunc_wire_205, {fourFunc_wire_207_0, fourFunc_wire_208_0});
xor_n #(2, 0, 0) XOR_67 (fourFunc_wire_187, {fourFunc_wire_209, fourFunc_wire_210_0});
xor_n #(2, 0, 0) XOR_68 (fourFunc_wire_209, {fourFunc_wire_211_0, fourFunc_wire_212_0});
xor_n #(2, 0, 0) XOR_69 (fourFunc_wire_213, {fourFunc_wire_214, fourFunc_wire_215});
xor_n #(2, 0, 0) XOR_70 (fourFunc_wire_214, {fourFunc_wire_216_0, fourFunc_wire_217});
xor_n #(2, 0, 0) XOR_71 (fourFunc_wire_195, {fourFunc_wire_218, fourFunc_wire_219_0});
xor_n #(2, 0, 0) XOR_72 (fourFunc_wire_218, {fourFunc_wire_220_0, fourFunc_wire_221_0});
xor_n #(2, 0, 0) XOR_73 (fourFunc_wire_199, {fourFunc_wire_222, fourFunc_wire_223_0});
xor_n #(2, 0, 0) XOR_74 (fourFunc_wire_222, {fourFunc_wire_224_0, fourFunc_wire_225_0});
xor_n #(2, 0, 0) XOR_75 (fourFunc_wire_203, {fourFunc_wire_226, fourFunc_wire_227_0});
xor_n #(2, 0, 0) XOR_76 (fourFunc_wire_226, {fourFunc_wire_228_0, fourFunc_wire_229_0});
xor_n #(2, 0, 0) XOR_77 (fourFunc_wire_207, {fourFunc_wire_230, fourFunc_wire_231_0});
xor_n #(2, 0, 0) XOR_78 (fourFunc_wire_230, {fourFunc_wire_232_0, fourFunc_wire_233_0});
xor_n #(2, 0, 0) XOR_79 (fourFunc_wire_211, {fourFunc_wire_234, fourFunc_wire_235_0});
xor_n #(2, 0, 0) XOR_80 (fourFunc_wire_234, {fourFunc_wire_236_0, fourFunc_wire_237_0});
xor_n #(2, 0, 0) XOR_81 (fourFunc_wire_216, {fourFunc_wire_238, fourFunc_wire_239_0});
xor_n #(2, 0, 0) XOR_82 (fourFunc_wire_238, {fourFunc_wire_240_0, fourFunc_wire_241_0});
xor_n #(2, 0, 0) XOR_83 (fourFunc_wire_242, {fourFunc_wire_243, fourFunc_wire_244});
xor_n #(2, 0, 0) XOR_84 (fourFunc_wire_243, {fourFunc_wire_245_0, fourFunc_wire_246});
xor_n #(2, 0, 0) XOR_85 (fourFunc_wire_224, {fourFunc_wire_247, fourFunc_wire_248_0});
xor_n #(2, 0, 0) XOR_86 (fourFunc_wire_247, {fourFunc_wire_249_0, fourFunc_wire_250_0});
xor_n #(2, 0, 0) XOR_87 (fourFunc_wire_228, {fourFunc_wire_251, fourFunc_wire_252_0});
xor_n #(2, 0, 0) XOR_88 (fourFunc_wire_251, {fourFunc_wire_253_0, fourFunc_wire_254_0});
xor_n #(2, 0, 0) XOR_89 (fourFunc_wire_232, {fourFunc_wire_255, fourFunc_wire_256_0});
xor_n #(2, 0, 0) XOR_90 (fourFunc_wire_255, {fourFunc_wire_257_0, fourFunc_wire_258_0});
xor_n #(2, 0, 0) XOR_91 (fourFunc_wire_236, {fourFunc_wire_259, fourFunc_wire_260_0});
xor_n #(2, 0, 0) XOR_92 (fourFunc_wire_259, {fourFunc_wire_261_0, fourFunc_wire_262_0});
xor_n #(2, 0, 0) XOR_93 (fourFunc_wire_240, {fourFunc_wire_263, fourFunc_wire_264_0});
xor_n #(2, 0, 0) XOR_94 (fourFunc_wire_263, {fourFunc_wire_265_0, fourFunc_wire_266_0});
xor_n #(2, 0, 0) XOR_95 (fourFunc_wire_245, {fourFunc_wire_267, fourFunc_wire_268_0});
xor_n #(2, 0, 0) XOR_96 (fourFunc_wire_267, {fourFunc_wire_269_0, fourFunc_wire_270_0});
xor_n #(2, 0, 0) XOR_97 (fourFunc_wire_271, {fourFunc_wire_272, fourFunc_wire_273});
xor_n #(2, 0, 0) XOR_98 (fourFunc_wire_272, {fourFunc_wire_274_0, fourFunc_wire_275});
xor_n #(2, 0, 0) XOR_99 (fourFunc_wire_253, {fourFunc_wire_276, fourFunc_wire_277_0});
xor_n #(2, 0, 0) XOR_100 (fourFunc_wire_276, {fourFunc_wire_278_0, fourFunc_wire_279_0});
xor_n #(2, 0, 0) XOR_101 (fourFunc_wire_257, {fourFunc_wire_280, fourFunc_wire_281_0});
xor_n #(2, 0, 0) XOR_102 (fourFunc_wire_280, {fourFunc_wire_122_0, fourFunc_wire_282_0});
xor_n #(2, 0, 0) XOR_103 (fourFunc_wire_261, {fourFunc_wire_283, fourFunc_wire_284_0});
xor_n #(2, 0, 0) XOR_104 (fourFunc_wire_283, {fourFunc_wire_285_0, fourFunc_wire_286_0});
xor_n #(2, 0, 0) XOR_105 (fourFunc_wire_265, {fourFunc_wire_287, fourFunc_wire_288_0});
xor_n #(2, 0, 0) XOR_106 (fourFunc_wire_287, {fourFunc_wire_289_0, fourFunc_wire_290_0});
xor_n #(2, 0, 0) XOR_107 (fourFunc_wire_269, {fourFunc_wire_291, fourFunc_wire_292_0});
xor_n #(2, 0, 0) XOR_108 (fourFunc_wire_291, {fourFunc_wire_293_0, fourFunc_wire_294_0});
xor_n #(2, 0, 0) XOR_109 (fourFunc_wire_274, {fourFunc_wire_295, fourFunc_wire_296_0});
xor_n #(2, 0, 0) XOR_110 (fourFunc_wire_295, {fourFunc_wire_297_0, fourFunc_wire_298_0});
xor_n #(2, 0, 0) XOR_111 (fourFunc_wire_299, {fourFunc_wire_300, fourFunc_wire_301});
xor_n #(2, 0, 0) XOR_112 (fourFunc_wire_300, {fourFunc_wire_302_0, fourFunc_wire_303});
xor_n #(2, 0, 0) XOR_113 (fourFunc_wire_285, {fourFunc_wire_304, fourFunc_wire_305_0});
xor_n #(2, 0, 0) XOR_114 (fourFunc_wire_304, {fourFunc_wire_306_0, fourFunc_wire_307_0});
xor_n #(2, 0, 0) XOR_115 (fourFunc_wire_289, {fourFunc_wire_308, fourFunc_wire_309_0});
xor_n #(2, 0, 0) XOR_116 (fourFunc_wire_308, {fourFunc_wire_310_0, fourFunc_wire_311_0});
xor_n #(2, 0, 0) XOR_117 (fourFunc_wire_293, {fourFunc_wire_312, fourFunc_wire_313_0});
xor_n #(2, 0, 0) XOR_118 (fourFunc_wire_312, {fourFunc_wire_314_0, fourFunc_wire_315_0});
xor_n #(2, 0, 0) XOR_119 (fourFunc_wire_297, {fourFunc_wire_316, fourFunc_wire_317_0});
xor_n #(2, 0, 0) XOR_120 (fourFunc_wire_316, {fourFunc_wire_318_0, fourFunc_wire_319_0});
xor_n #(2, 0, 0) XOR_121 (fourFunc_wire_302, {fourFunc_wire_320, fourFunc_wire_321_0});
xor_n #(2, 0, 0) XOR_122 (fourFunc_wire_320, {fourFunc_wire_322_0, fourFunc_wire_323_0});
xor_n #(2, 0, 0) XOR_123 (fourFunc_wire_324, {fourFunc_wire_325, fourFunc_wire_326});
xor_n #(2, 0, 0) XOR_124 (fourFunc_wire_325, {fourFunc_wire_327_0, fourFunc_wire_328_0});
and_n #(2, 0, 0) AND_14 (fourFunc_wire_121, {fourFunc_wire_54_2, fourFunc_wire_53_2});
and_n #(2, 0, 0) AND_15 (fourFunc_wire_329, {fourFunc_wire_121_1, fourFunc_wire_330});
and_n #(2, 0, 0) AND_16 (fourFunc_wire_100, {fourFunc_wire_98_1, fourFunc_wire_59_2});
or_n #(2, 0, 0) OR_9 (fourFunc_wire_118, {fourFunc_wire_331, fourFunc_wire_329});
and_n #(2, 0, 0) AND_17 (fourFunc_wire_332, {fourFunc_wire_118_1, fourFunc_wire_333});
and_n #(2, 0, 0) AND_18 (fourFunc_wire_331, {fourFunc_wire_94_2, fourFunc_wire_95_2});
or_n #(2, 0, 0) OR_10 (fourFunc_wire_330, {fourFunc_wire_94_3, fourFunc_wire_95_3});
or_n #(2, 0, 0) OR_11 (fourFunc_wire_115, {fourFunc_wire_334, fourFunc_wire_332});
and_n #(2, 0, 0) AND_19 (fourFunc_wire_335, {fourFunc_wire_115_1, fourFunc_wire_336});
and_n #(2, 0, 0) AND_20 (fourFunc_wire_334, {fourFunc_wire_89_2, fourFunc_wire_90_2});
or_n #(2, 0, 0) OR_12 (fourFunc_wire_333, {fourFunc_wire_89_3, fourFunc_wire_90_3});
or_n #(2, 0, 0) OR_13 (fourFunc_wire_112, {fourFunc_wire_337, fourFunc_wire_335});
and_n #(2, 0, 0) AND_21 (fourFunc_wire_338, {fourFunc_wire_112_1, fourFunc_wire_339});
and_n #(2, 0, 0) AND_22 (fourFunc_wire_337, {fourFunc_wire_84_2, fourFunc_wire_85_2});
or_n #(2, 0, 0) OR_14 (fourFunc_wire_336, {fourFunc_wire_84_3, fourFunc_wire_85_3});
or_n #(2, 0, 0) OR_15 (fourFunc_wire_109, {fourFunc_wire_340, fourFunc_wire_338});
and_n #(2, 0, 0) AND_23 (fourFunc_wire_341, {fourFunc_wire_109_1, fourFunc_wire_342});
and_n #(2, 0, 0) AND_24 (fourFunc_wire_340, {fourFunc_wire_79_2, fourFunc_wire_80_2});
or_n #(2, 0, 0) OR_16 (fourFunc_wire_339, {fourFunc_wire_79_3, fourFunc_wire_80_3});
or_n #(2, 0, 0) OR_17 (fourFunc_wire_106, {fourFunc_wire_343, fourFunc_wire_341});
and_n #(2, 0, 0) AND_25 (fourFunc_wire_344, {fourFunc_wire_106_1, fourFunc_wire_345});
and_n #(2, 0, 0) AND_26 (fourFunc_wire_343, {fourFunc_wire_74_2, fourFunc_wire_75_2});
or_n #(2, 0, 0) OR_18 (fourFunc_wire_342, {fourFunc_wire_74_3, fourFunc_wire_75_3});
or_n #(2, 0, 0) OR_19 (fourFunc_wire_103, {fourFunc_wire_346, fourFunc_wire_344});
and_n #(2, 0, 0) AND_27 (fourFunc_wire_347, {fourFunc_wire_103_1, fourFunc_wire_348});
and_n #(2, 0, 0) AND_28 (fourFunc_wire_346, {fourFunc_wire_69_2, fourFunc_wire_70_2});
or_n #(2, 0, 0) OR_20 (fourFunc_wire_345, {fourFunc_wire_69_3, fourFunc_wire_70_3});
or_n #(2, 0, 0) OR_21 (fourFunc_wire_98, {fourFunc_wire_349, fourFunc_wire_347});
and_n #(2, 0, 0) AND_29 (fourFunc_wire_349, {fourFunc_wire_64_2, fourFunc_wire_65_2});
or_n #(2, 0, 0) OR_22 (fourFunc_wire_348, {fourFunc_wire_64_3, fourFunc_wire_65_3});
and_n #(3, 0, 0) AND_30 (fourFunc_wire_301, {fourFunc_wire_324_0, fourFunc_wire_350_0, fourFunc_wire_53_3});
and_n #(2, 0, 0) AND_31 (fourFunc_wire_351, {fourFunc_wire_324_1, fourFunc_wire_53_4});
and_n #(2, 0, 0) AND_32 (fourFunc_wire_352, {fourFunc_wire_302_1, fourFunc_wire_95_4});
or_n #(2, 0, 0) OR_23 (fourFunc_wire_353, {fourFunc_wire_302_2, fourFunc_wire_95_5});
and_n #(2, 0, 0) AND_33 (fourFunc_wire_354, {fourFunc_wire_297_1, fourFunc_wire_296_1});
or_n #(2, 0, 0) OR_24 (fourFunc_wire_355, {fourFunc_wire_297_2, fourFunc_wire_296_2});
and_n #(2, 0, 0) AND_34 (fourFunc_wire_356, {fourFunc_wire_293_1, fourFunc_wire_292_1});
or_n #(2, 0, 0) OR_25 (fourFunc_wire_357, {fourFunc_wire_293_2, fourFunc_wire_292_2});
and_n #(2, 0, 0) AND_35 (fourFunc_wire_358, {fourFunc_wire_289_1, fourFunc_wire_288_1});
or_n #(2, 0, 0) OR_26 (fourFunc_wire_359, {fourFunc_wire_289_2, fourFunc_wire_288_2});
and_n #(2, 0, 0) AND_36 (fourFunc_wire_360, {fourFunc_wire_285_1, fourFunc_wire_284_1});
or_n #(2, 0, 0) OR_27 (fourFunc_wire_361, {fourFunc_wire_285_2, fourFunc_wire_284_2});
and_n #(2, 0, 0) AND_37 (fourFunc_wire_362, {fourFunc_wire_122_1, fourFunc_wire_281_1});
or_n #(2, 0, 0) OR_28 (fourFunc_wire_363, {fourFunc_wire_122_2, fourFunc_wire_281_2});
and_n #(3, 0, 0) AND_38 (fourFunc_wire_273, {fourFunc_wire_299_0, fourFunc_wire_364_0, fourFunc_wire_53_5});
and_n #(2, 0, 0) AND_39 (fourFunc_wire_365, {fourFunc_wire_299_1, fourFunc_wire_53_6});
and_n #(2, 0, 0) AND_40 (fourFunc_wire_366, {fourFunc_wire_274_1, fourFunc_wire_95_6});
or_n #(2, 0, 0) OR_29 (fourFunc_wire_367, {fourFunc_wire_274_2, fourFunc_wire_95_7});
and_n #(2, 0, 0) AND_41 (fourFunc_wire_368, {fourFunc_wire_269_1, fourFunc_wire_268_1});
or_n #(2, 0, 0) OR_30 (fourFunc_wire_369, {fourFunc_wire_269_2, fourFunc_wire_268_2});
and_n #(2, 0, 0) AND_42 (fourFunc_wire_370, {fourFunc_wire_265_1, fourFunc_wire_264_1});
or_n #(2, 0, 0) OR_31 (fourFunc_wire_371, {fourFunc_wire_265_2, fourFunc_wire_264_2});
and_n #(2, 0, 0) AND_43 (fourFunc_wire_372, {fourFunc_wire_261_1, fourFunc_wire_260_1});
or_n #(2, 0, 0) OR_32 (fourFunc_wire_373, {fourFunc_wire_261_2, fourFunc_wire_260_2});
and_n #(2, 0, 0) AND_44 (fourFunc_wire_374, {fourFunc_wire_257_1, fourFunc_wire_256_1});
or_n #(2, 0, 0) OR_33 (fourFunc_wire_375, {fourFunc_wire_257_2, fourFunc_wire_256_2});
and_n #(2, 0, 0) AND_45 (fourFunc_wire_376, {fourFunc_wire_253_1, fourFunc_wire_252_1});
or_n #(2, 0, 0) OR_34 (fourFunc_wire_377, {fourFunc_wire_253_2, fourFunc_wire_252_2});
and_n #(3, 0, 0) AND_46 (fourFunc_wire_244, {fourFunc_wire_271_0, fourFunc_wire_378_0, fourFunc_wire_53_7});
and_n #(2, 0, 0) AND_47 (fourFunc_wire_379, {fourFunc_wire_271_1, fourFunc_wire_53_8});
and_n #(2, 0, 0) AND_48 (fourFunc_wire_380, {fourFunc_wire_245_1, fourFunc_wire_95_8});
or_n #(2, 0, 0) OR_35 (fourFunc_wire_381, {fourFunc_wire_245_2, fourFunc_wire_95_9});
and_n #(2, 0, 0) AND_49 (fourFunc_wire_382, {fourFunc_wire_240_1, fourFunc_wire_239_1});
or_n #(2, 0, 0) OR_36 (fourFunc_wire_383, {fourFunc_wire_240_2, fourFunc_wire_239_2});
and_n #(2, 0, 0) AND_50 (fourFunc_wire_384, {fourFunc_wire_236_1, fourFunc_wire_235_1});
or_n #(2, 0, 0) OR_37 (fourFunc_wire_385, {fourFunc_wire_236_2, fourFunc_wire_235_2});
and_n #(2, 0, 0) AND_51 (fourFunc_wire_386, {fourFunc_wire_232_1, fourFunc_wire_231_1});
or_n #(2, 0, 0) OR_38 (fourFunc_wire_387, {fourFunc_wire_232_2, fourFunc_wire_231_2});
and_n #(2, 0, 0) AND_52 (fourFunc_wire_388, {fourFunc_wire_228_1, fourFunc_wire_227_1});
or_n #(2, 0, 0) OR_39 (fourFunc_wire_389, {fourFunc_wire_228_2, fourFunc_wire_227_2});
and_n #(2, 0, 0) AND_53 (fourFunc_wire_390, {fourFunc_wire_224_1, fourFunc_wire_223_1});
or_n #(2, 0, 0) OR_40 (fourFunc_wire_391, {fourFunc_wire_224_2, fourFunc_wire_223_2});
and_n #(3, 0, 0) AND_54 (fourFunc_wire_215, {fourFunc_wire_242_0, fourFunc_wire_392_0, fourFunc_wire_53_9});
and_n #(2, 0, 0) AND_55 (fourFunc_wire_393, {fourFunc_wire_242_1, fourFunc_wire_53_10});
and_n #(2, 0, 0) AND_56 (fourFunc_wire_394, {fourFunc_wire_216_1, fourFunc_wire_95_10});
or_n #(2, 0, 0) OR_41 (fourFunc_wire_395, {fourFunc_wire_216_2, fourFunc_wire_95_11});
and_n #(2, 0, 0) AND_57 (fourFunc_wire_396, {fourFunc_wire_211_1, fourFunc_wire_210_1});
or_n #(2, 0, 0) OR_42 (fourFunc_wire_397, {fourFunc_wire_211_2, fourFunc_wire_210_2});
and_n #(2, 0, 0) AND_58 (fourFunc_wire_398, {fourFunc_wire_207_1, fourFunc_wire_206_1});
or_n #(2, 0, 0) OR_43 (fourFunc_wire_399, {fourFunc_wire_207_2, fourFunc_wire_206_2});
and_n #(2, 0, 0) AND_59 (fourFunc_wire_400, {fourFunc_wire_203_1, fourFunc_wire_202_1});
or_n #(2, 0, 0) OR_44 (fourFunc_wire_401, {fourFunc_wire_203_2, fourFunc_wire_202_2});
and_n #(2, 0, 0) AND_60 (fourFunc_wire_402, {fourFunc_wire_199_1, fourFunc_wire_198_1});
or_n #(2, 0, 0) OR_45 (fourFunc_wire_403, {fourFunc_wire_199_2, fourFunc_wire_198_2});
and_n #(2, 0, 0) AND_61 (fourFunc_wire_404, {fourFunc_wire_195_1, fourFunc_wire_194_1});
or_n #(2, 0, 0) OR_46 (fourFunc_wire_405, {fourFunc_wire_195_2, fourFunc_wire_194_2});
and_n #(3, 0, 0) AND_62 (fourFunc_wire_186, {fourFunc_wire_213_0, fourFunc_wire_406_0, fourFunc_wire_53_11});
and_n #(2, 0, 0) AND_63 (fourFunc_wire_407, {fourFunc_wire_213_1, fourFunc_wire_53_12});
and_n #(2, 0, 0) AND_64 (fourFunc_wire_408, {fourFunc_wire_187_1, fourFunc_wire_95_12});
or_n #(2, 0, 0) OR_47 (fourFunc_wire_409, {fourFunc_wire_187_2, fourFunc_wire_95_13});
and_n #(2, 0, 0) AND_65 (fourFunc_wire_410, {fourFunc_wire_182_1, fourFunc_wire_181_1});
or_n #(2, 0, 0) OR_48 (fourFunc_wire_411, {fourFunc_wire_182_2, fourFunc_wire_181_2});
and_n #(2, 0, 0) AND_66 (fourFunc_wire_412, {fourFunc_wire_178_1, fourFunc_wire_177_1});
or_n #(2, 0, 0) OR_49 (fourFunc_wire_413, {fourFunc_wire_178_2, fourFunc_wire_177_2});
and_n #(2, 0, 0) AND_67 (fourFunc_wire_414, {fourFunc_wire_174_1, fourFunc_wire_173_1});
or_n #(2, 0, 0) OR_50 (fourFunc_wire_415, {fourFunc_wire_174_2, fourFunc_wire_173_2});
and_n #(2, 0, 0) AND_68 (fourFunc_wire_416, {fourFunc_wire_170_1, fourFunc_wire_169_1});
or_n #(2, 0, 0) OR_51 (fourFunc_wire_417, {fourFunc_wire_170_2, fourFunc_wire_169_2});
and_n #(2, 0, 0) AND_69 (fourFunc_wire_418, {fourFunc_wire_166_1, fourFunc_wire_165_1});
or_n #(2, 0, 0) OR_52 (fourFunc_wire_419, {fourFunc_wire_166_2, fourFunc_wire_165_2});
and_n #(3, 0, 0) AND_70 (fourFunc_wire_157, {fourFunc_wire_184_0, fourFunc_wire_420_0, fourFunc_wire_53_13});
and_n #(2, 0, 0) AND_71 (fourFunc_wire_421, {fourFunc_wire_184_1, fourFunc_wire_53_14});
and_n #(2, 0, 0) AND_72 (fourFunc_wire_422, {fourFunc_wire_158_1, fourFunc_wire_95_14});
or_n #(2, 0, 0) OR_53 (fourFunc_wire_423, {fourFunc_wire_158_2, fourFunc_wire_95_15});
and_n #(2, 0, 0) AND_73 (fourFunc_wire_424, {fourFunc_wire_153_1, fourFunc_wire_152_1});
or_n #(2, 0, 0) OR_54 (fourFunc_wire_425, {fourFunc_wire_153_2, fourFunc_wire_152_2});
and_n #(2, 0, 0) AND_74 (fourFunc_wire_426, {fourFunc_wire_148_1, fourFunc_wire_147_1});
or_n #(2, 0, 0) OR_55 (fourFunc_wire_427, {fourFunc_wire_148_2, fourFunc_wire_147_2});
and_n #(2, 0, 0) AND_75 (fourFunc_wire_428, {fourFunc_wire_143_1, fourFunc_wire_142_1});
or_n #(2, 0, 0) OR_56 (fourFunc_wire_429, {fourFunc_wire_143_2, fourFunc_wire_142_2});
and_n #(2, 0, 0) AND_76 (fourFunc_wire_430, {fourFunc_wire_138_1, fourFunc_wire_137_1});
or_n #(2, 0, 0) OR_57 (fourFunc_wire_431, {fourFunc_wire_138_2, fourFunc_wire_137_2});
and_n #(2, 0, 0) AND_77 (fourFunc_wire_432, {fourFunc_wire_133_1, fourFunc_wire_132_1});
or_n #(2, 0, 0) OR_58 (fourFunc_wire_433, {fourFunc_wire_133_2, fourFunc_wire_132_2});
and_n #(2, 0, 0) AND_78 (fourFunc_wire_306, {fourFunc_wire_434_0, fourFunc_wire_65_4});
and_n #(2, 0, 0) AND_79 (fourFunc_wire_435, {fourFunc_wire_306_1, fourFunc_wire_436});
and_n #(2, 0, 0) AND_80 (fourFunc_wire_310, {fourFunc_wire_434_1, fourFunc_wire_70_4});
and_n #(2, 0, 0) AND_81 (fourFunc_wire_437, {fourFunc_wire_310_1, fourFunc_wire_438});
and_n #(2, 0, 0) AND_82 (fourFunc_wire_314, {fourFunc_wire_434_2, fourFunc_wire_75_4});
and_n #(2, 0, 0) AND_83 (fourFunc_wire_439, {fourFunc_wire_314_1, fourFunc_wire_440});
and_n #(2, 0, 0) AND_84 (fourFunc_wire_318, {fourFunc_wire_434_3, fourFunc_wire_80_4});
and_n #(2, 0, 0) AND_85 (fourFunc_wire_441, {fourFunc_wire_318_1, fourFunc_wire_442});
and_n #(2, 0, 0) AND_86 (fourFunc_wire_322, {fourFunc_wire_434_4, fourFunc_wire_85_4});
and_n #(2, 0, 0) AND_87 (fourFunc_wire_443, {fourFunc_wire_322_1, fourFunc_wire_444});
and_n #(2, 0, 0) AND_88 (fourFunc_wire_327, {fourFunc_wire_434_5, fourFunc_wire_90_4});
and_n #(2, 0, 0) AND_89 (fourFunc_wire_445, {fourFunc_wire_327_1, fourFunc_wire_328_1});
and_n #(2, 0, 0) AND_90 (fourFunc_wire_278, {fourFunc_wire_124_1, fourFunc_wire_123_1});
and_n #(2, 0, 0) AND_91 (fourFunc_wire_124, {fourFunc_wire_446_0, fourFunc_wire_65_5});
and_n #(2, 0, 0) AND_92 (fourFunc_wire_307, {fourFunc_wire_446_1, fourFunc_wire_70_5});
and_n #(2, 0, 0) AND_93 (fourFunc_wire_447, {fourFunc_wire_307_1, fourFunc_wire_305_1});
or_n #(2, 0, 0) OR_59 (fourFunc_wire_436, {fourFunc_wire_307_2, fourFunc_wire_305_2});
and_n #(2, 0, 0) AND_94 (fourFunc_wire_311, {fourFunc_wire_446_2, fourFunc_wire_75_5});
and_n #(2, 0, 0) AND_95 (fourFunc_wire_448, {fourFunc_wire_311_1, fourFunc_wire_309_1});
or_n #(2, 0, 0) OR_60 (fourFunc_wire_438, {fourFunc_wire_311_2, fourFunc_wire_309_2});
and_n #(2, 0, 0) AND_96 (fourFunc_wire_315, {fourFunc_wire_446_3, fourFunc_wire_80_5});
and_n #(2, 0, 0) AND_97 (fourFunc_wire_449, {fourFunc_wire_315_1, fourFunc_wire_313_1});
or_n #(2, 0, 0) OR_61 (fourFunc_wire_440, {fourFunc_wire_315_2, fourFunc_wire_313_2});
and_n #(2, 0, 0) AND_98 (fourFunc_wire_319, {fourFunc_wire_446_4, fourFunc_wire_85_5});
and_n #(2, 0, 0) AND_99 (fourFunc_wire_450, {fourFunc_wire_319_1, fourFunc_wire_317_1});
or_n #(2, 0, 0) OR_62 (fourFunc_wire_442, {fourFunc_wire_319_2, fourFunc_wire_317_2});
and_n #(2, 0, 0) AND_100 (fourFunc_wire_323, {fourFunc_wire_446_5, fourFunc_wire_90_5});
and_n #(2, 0, 0) AND_101 (fourFunc_wire_451, {fourFunc_wire_323_1, fourFunc_wire_321_1});
or_n #(2, 0, 0) OR_63 (fourFunc_wire_444, {fourFunc_wire_323_2, fourFunc_wire_321_2});
and_n #(2, 0, 0) AND_102 (fourFunc_wire_328, {fourFunc_wire_446_6, fourFunc_wire_95_16});
and_n #(4, 0, 0) AND_103 (fourFunc_wire_326, {fourFunc_wire_434_6, fourFunc_wire_446_7, fourFunc_wire_53_15, fourFunc_wire_95_17});
and_n #(2, 0, 0) AND_104 (fourFunc_wire_279, {fourFunc_wire_350_1, fourFunc_wire_65_6});
and_n #(2, 0, 0) AND_105 (fourFunc_wire_452, {fourFunc_wire_279_1, fourFunc_wire_453});
and_n #(2, 0, 0) AND_106 (fourFunc_wire_282, {fourFunc_wire_350_2, fourFunc_wire_70_6});
and_n #(2, 0, 0) AND_107 (fourFunc_wire_454, {fourFunc_wire_282_1, fourFunc_wire_363});
and_n #(2, 0, 0) AND_108 (fourFunc_wire_286, {fourFunc_wire_350_3, fourFunc_wire_75_6});
and_n #(2, 0, 0) AND_109 (fourFunc_wire_455, {fourFunc_wire_286_1, fourFunc_wire_361});
and_n #(2, 0, 0) AND_110 (fourFunc_wire_290, {fourFunc_wire_350_4, fourFunc_wire_80_6});
and_n #(2, 0, 0) AND_111 (fourFunc_wire_456, {fourFunc_wire_290_1, fourFunc_wire_359});
and_n #(2, 0, 0) AND_112 (fourFunc_wire_294, {fourFunc_wire_350_5, fourFunc_wire_85_6});
and_n #(2, 0, 0) AND_113 (fourFunc_wire_457, {fourFunc_wire_294_1, fourFunc_wire_357});
and_n #(2, 0, 0) AND_114 (fourFunc_wire_298, {fourFunc_wire_350_6, fourFunc_wire_90_6});
and_n #(2, 0, 0) AND_115 (fourFunc_wire_458, {fourFunc_wire_298_1, fourFunc_wire_355});
and_n #(2, 0, 0) AND_116 (fourFunc_wire_303, {fourFunc_wire_350_7, fourFunc_wire_95_18});
and_n #(2, 0, 0) AND_117 (fourFunc_wire_250, {fourFunc_wire_364_1, fourFunc_wire_65_7});
and_n #(2, 0, 0) AND_118 (fourFunc_wire_459, {fourFunc_wire_250_1, fourFunc_wire_460});
and_n #(2, 0, 0) AND_119 (fourFunc_wire_254, {fourFunc_wire_364_2, fourFunc_wire_70_7});
and_n #(2, 0, 0) AND_120 (fourFunc_wire_461, {fourFunc_wire_254_1, fourFunc_wire_377});
and_n #(2, 0, 0) AND_121 (fourFunc_wire_258, {fourFunc_wire_364_3, fourFunc_wire_75_7});
and_n #(2, 0, 0) AND_122 (fourFunc_wire_462, {fourFunc_wire_258_1, fourFunc_wire_375});
and_n #(2, 0, 0) AND_123 (fourFunc_wire_262, {fourFunc_wire_364_4, fourFunc_wire_80_7});
and_n #(2, 0, 0) AND_124 (fourFunc_wire_463, {fourFunc_wire_262_1, fourFunc_wire_373});
and_n #(2, 0, 0) AND_125 (fourFunc_wire_266, {fourFunc_wire_364_5, fourFunc_wire_85_7});
and_n #(2, 0, 0) AND_126 (fourFunc_wire_464, {fourFunc_wire_266_1, fourFunc_wire_371});
and_n #(2, 0, 0) AND_127 (fourFunc_wire_270, {fourFunc_wire_364_6, fourFunc_wire_90_7});
and_n #(2, 0, 0) AND_128 (fourFunc_wire_465, {fourFunc_wire_270_1, fourFunc_wire_369});
and_n #(2, 0, 0) AND_129 (fourFunc_wire_275, {fourFunc_wire_364_7, fourFunc_wire_95_19});
and_n #(2, 0, 0) AND_130 (fourFunc_wire_221, {fourFunc_wire_378_1, fourFunc_wire_65_8});
and_n #(2, 0, 0) AND_131 (fourFunc_wire_466, {fourFunc_wire_221_1, fourFunc_wire_467});
and_n #(2, 0, 0) AND_132 (fourFunc_wire_225, {fourFunc_wire_378_2, fourFunc_wire_70_8});
and_n #(2, 0, 0) AND_133 (fourFunc_wire_468, {fourFunc_wire_225_1, fourFunc_wire_391});
and_n #(2, 0, 0) AND_134 (fourFunc_wire_229, {fourFunc_wire_378_3, fourFunc_wire_75_8});
and_n #(2, 0, 0) AND_135 (fourFunc_wire_469, {fourFunc_wire_229_1, fourFunc_wire_389});
and_n #(2, 0, 0) AND_136 (fourFunc_wire_233, {fourFunc_wire_378_4, fourFunc_wire_80_8});
and_n #(2, 0, 0) AND_137 (fourFunc_wire_470, {fourFunc_wire_233_1, fourFunc_wire_387});
and_n #(2, 0, 0) AND_138 (fourFunc_wire_237, {fourFunc_wire_378_5, fourFunc_wire_85_8});
and_n #(2, 0, 0) AND_139 (fourFunc_wire_471, {fourFunc_wire_237_1, fourFunc_wire_385});
and_n #(2, 0, 0) AND_140 (fourFunc_wire_241, {fourFunc_wire_378_6, fourFunc_wire_90_8});
and_n #(2, 0, 0) AND_141 (fourFunc_wire_472, {fourFunc_wire_241_1, fourFunc_wire_383});
and_n #(2, 0, 0) AND_142 (fourFunc_wire_246, {fourFunc_wire_378_7, fourFunc_wire_95_20});
and_n #(2, 0, 0) AND_143 (fourFunc_wire_192, {fourFunc_wire_392_1, fourFunc_wire_65_9});
and_n #(2, 0, 0) AND_144 (fourFunc_wire_473, {fourFunc_wire_192_1, fourFunc_wire_474});
and_n #(2, 0, 0) AND_145 (fourFunc_wire_196, {fourFunc_wire_392_2, fourFunc_wire_70_9});
and_n #(2, 0, 0) AND_146 (fourFunc_wire_475, {fourFunc_wire_196_1, fourFunc_wire_405});
and_n #(2, 0, 0) AND_147 (fourFunc_wire_200, {fourFunc_wire_392_3, fourFunc_wire_75_9});
and_n #(2, 0, 0) AND_148 (fourFunc_wire_476, {fourFunc_wire_200_1, fourFunc_wire_403});
and_n #(2, 0, 0) AND_149 (fourFunc_wire_204, {fourFunc_wire_392_4, fourFunc_wire_80_9});
and_n #(2, 0, 0) AND_150 (fourFunc_wire_477, {fourFunc_wire_204_1, fourFunc_wire_401});
and_n #(2, 0, 0) AND_151 (fourFunc_wire_208, {fourFunc_wire_392_5, fourFunc_wire_85_9});
and_n #(2, 0, 0) AND_152 (fourFunc_wire_478, {fourFunc_wire_208_1, fourFunc_wire_399});
and_n #(2, 0, 0) AND_153 (fourFunc_wire_212, {fourFunc_wire_392_6, fourFunc_wire_90_9});
and_n #(2, 0, 0) AND_154 (fourFunc_wire_479, {fourFunc_wire_212_1, fourFunc_wire_397});
and_n #(2, 0, 0) AND_155 (fourFunc_wire_217, {fourFunc_wire_392_7, fourFunc_wire_95_21});
and_n #(2, 0, 0) AND_156 (fourFunc_wire_163, {fourFunc_wire_406_1, fourFunc_wire_65_10});
and_n #(2, 0, 0) AND_157 (fourFunc_wire_480, {fourFunc_wire_163_1, fourFunc_wire_481});
and_n #(2, 0, 0) AND_158 (fourFunc_wire_167, {fourFunc_wire_406_2, fourFunc_wire_70_10});
and_n #(2, 0, 0) AND_159 (fourFunc_wire_482, {fourFunc_wire_167_1, fourFunc_wire_419});
and_n #(2, 0, 0) AND_160 (fourFunc_wire_171, {fourFunc_wire_406_3, fourFunc_wire_75_10});
and_n #(2, 0, 0) AND_161 (fourFunc_wire_483, {fourFunc_wire_171_1, fourFunc_wire_417});
and_n #(2, 0, 0) AND_162 (fourFunc_wire_175, {fourFunc_wire_406_4, fourFunc_wire_80_10});
and_n #(2, 0, 0) AND_163 (fourFunc_wire_484, {fourFunc_wire_175_1, fourFunc_wire_415});
and_n #(2, 0, 0) AND_164 (fourFunc_wire_179, {fourFunc_wire_406_5, fourFunc_wire_85_10});
and_n #(2, 0, 0) AND_165 (fourFunc_wire_485, {fourFunc_wire_179_1, fourFunc_wire_413});
and_n #(2, 0, 0) AND_166 (fourFunc_wire_183, {fourFunc_wire_406_6, fourFunc_wire_90_10});
and_n #(2, 0, 0) AND_167 (fourFunc_wire_486, {fourFunc_wire_183_1, fourFunc_wire_411});
and_n #(2, 0, 0) AND_168 (fourFunc_wire_188, {fourFunc_wire_406_7, fourFunc_wire_95_22});
and_n #(2, 0, 0) AND_169 (fourFunc_wire_129, {fourFunc_wire_420_1, fourFunc_wire_65_11});
and_n #(2, 0, 0) AND_170 (fourFunc_wire_487, {fourFunc_wire_129_1, fourFunc_wire_488});
and_n #(2, 0, 0) AND_171 (fourFunc_wire_134, {fourFunc_wire_420_2, fourFunc_wire_70_11});
and_n #(2, 0, 0) AND_172 (fourFunc_wire_489, {fourFunc_wire_134_1, fourFunc_wire_433});
and_n #(2, 0, 0) AND_173 (fourFunc_wire_139, {fourFunc_wire_420_3, fourFunc_wire_75_11});
and_n #(2, 0, 0) AND_174 (fourFunc_wire_490, {fourFunc_wire_139_1, fourFunc_wire_431});
and_n #(2, 0, 0) AND_175 (fourFunc_wire_144, {fourFunc_wire_420_4, fourFunc_wire_80_11});
and_n #(2, 0, 0) AND_176 (fourFunc_wire_491, {fourFunc_wire_144_1, fourFunc_wire_429});
and_n #(2, 0, 0) AND_177 (fourFunc_wire_149, {fourFunc_wire_420_5, fourFunc_wire_85_11});
and_n #(2, 0, 0) AND_178 (fourFunc_wire_492, {fourFunc_wire_149_1, fourFunc_wire_427});
and_n #(2, 0, 0) AND_179 (fourFunc_wire_154, {fourFunc_wire_420_6, fourFunc_wire_90_11});
and_n #(2, 0, 0) AND_180 (fourFunc_wire_493, {fourFunc_wire_154_1, fourFunc_wire_425});
and_n #(2, 0, 0) AND_181 (fourFunc_wire_159, {fourFunc_wire_420_7, fourFunc_wire_95_23});
and_n #(2, 0, 0) AND_182 (fourFunc_wire_494, {fourFunc_wire_278_1, fourFunc_wire_277_1});
or_n #(2, 0, 0) OR_64 (fourFunc_wire_453, {fourFunc_wire_278_2, fourFunc_wire_277_2});
or_n #(2, 0, 0) OR_65 (fourFunc_wire_249, {fourFunc_wire_494, fourFunc_wire_452});
and_n #(2, 0, 0) AND_183 (fourFunc_wire_495, {fourFunc_wire_249_1, fourFunc_wire_248_1});
or_n #(2, 0, 0) OR_66 (fourFunc_wire_460, {fourFunc_wire_249_2, fourFunc_wire_248_2});
or_n #(2, 0, 0) OR_67 (fourFunc_wire_220, {fourFunc_wire_495, fourFunc_wire_459});
and_n #(2, 0, 0) AND_184 (fourFunc_wire_496, {fourFunc_wire_220_1, fourFunc_wire_219_1});
or_n #(2, 0, 0) OR_68 (fourFunc_wire_467, {fourFunc_wire_220_2, fourFunc_wire_219_2});
or_n #(2, 0, 0) OR_69 (fourFunc_wire_191, {fourFunc_wire_496, fourFunc_wire_466});
and_n #(2, 0, 0) AND_185 (fourFunc_wire_497, {fourFunc_wire_191_1, fourFunc_wire_190_1});
or_n #(2, 0, 0) OR_70 (fourFunc_wire_474, {fourFunc_wire_191_2, fourFunc_wire_190_2});
or_n #(2, 0, 0) OR_71 (fourFunc_wire_162, {fourFunc_wire_497, fourFunc_wire_473});
and_n #(2, 0, 0) AND_186 (fourFunc_wire_498, {fourFunc_wire_162_1, fourFunc_wire_161_1});
or_n #(2, 0, 0) OR_72 (fourFunc_wire_481, {fourFunc_wire_162_2, fourFunc_wire_161_2});
or_n #(2, 0, 0) OR_73 (fourFunc_wire_128, {fourFunc_wire_498, fourFunc_wire_480});
and_n #(2, 0, 0) AND_187 (fourFunc_wire_499, {fourFunc_wire_128_1, fourFunc_wire_127_1});
or_n #(2, 0, 0) OR_74 (fourFunc_wire_488, {fourFunc_wire_128_2, fourFunc_wire_127_2});
or_n #(2, 0, 0) OR_75 (fourFunc_wire_321, {fourFunc_wire_445, fourFunc_wire_500});
and_n #(4, 0, 0) AND_188 (fourFunc_wire_500, {fourFunc_wire_434_7, fourFunc_wire_446_8, fourFunc_wire_53_16, fourFunc_wire_95_24});
or_n #(2, 0, 0) OR_76 (fourFunc_wire_317, {fourFunc_wire_451, fourFunc_wire_443});
or_n #(2, 0, 0) OR_77 (fourFunc_wire_313, {fourFunc_wire_450, fourFunc_wire_441});
or_n #(2, 0, 0) OR_78 (fourFunc_wire_309, {fourFunc_wire_449, fourFunc_wire_439});
or_n #(2, 0, 0) OR_79 (fourFunc_wire_305, {fourFunc_wire_448, fourFunc_wire_437});
or_n #(2, 0, 0) OR_80 (fourFunc_wire_123, {fourFunc_wire_447, fourFunc_wire_435});
and_n #(2, 0, 0) AND_189 (fourFunc_wire_296, {fourFunc_wire_501, fourFunc_wire_350_8});
or_n #(2, 0, 0) OR_81 (fourFunc_wire_501, {fourFunc_wire_352, fourFunc_wire_502});
and_n #(2, 0, 0) AND_190 (fourFunc_wire_502, {fourFunc_wire_351, fourFunc_wire_353});
or_n #(2, 0, 0) OR_82 (fourFunc_wire_292, {fourFunc_wire_354, fourFunc_wire_458});
or_n #(2, 0, 0) OR_83 (fourFunc_wire_288, {fourFunc_wire_356, fourFunc_wire_457});
or_n #(2, 0, 0) OR_84 (fourFunc_wire_284, {fourFunc_wire_358, fourFunc_wire_456});
or_n #(2, 0, 0) OR_85 (fourFunc_wire_281, {fourFunc_wire_360, fourFunc_wire_455});
or_n #(2, 0, 0) OR_86 (fourFunc_wire_277, {fourFunc_wire_362, fourFunc_wire_454});
and_n #(2, 0, 0) AND_191 (fourFunc_wire_268, {fourFunc_wire_503, fourFunc_wire_364_8});
or_n #(2, 0, 0) OR_87 (fourFunc_wire_503, {fourFunc_wire_366, fourFunc_wire_504});
and_n #(2, 0, 0) AND_192 (fourFunc_wire_504, {fourFunc_wire_365, fourFunc_wire_367});
or_n #(2, 0, 0) OR_88 (fourFunc_wire_264, {fourFunc_wire_368, fourFunc_wire_465});
or_n #(2, 0, 0) OR_89 (fourFunc_wire_260, {fourFunc_wire_370, fourFunc_wire_464});
or_n #(2, 0, 0) OR_90 (fourFunc_wire_256, {fourFunc_wire_372, fourFunc_wire_463});
or_n #(2, 0, 0) OR_91 (fourFunc_wire_252, {fourFunc_wire_374, fourFunc_wire_462});
or_n #(2, 0, 0) OR_92 (fourFunc_wire_248, {fourFunc_wire_376, fourFunc_wire_461});
and_n #(2, 0, 0) AND_193 (fourFunc_wire_239, {fourFunc_wire_505, fourFunc_wire_378_8});
or_n #(2, 0, 0) OR_93 (fourFunc_wire_505, {fourFunc_wire_380, fourFunc_wire_506});
and_n #(2, 0, 0) AND_194 (fourFunc_wire_506, {fourFunc_wire_379, fourFunc_wire_381});
or_n #(2, 0, 0) OR_94 (fourFunc_wire_235, {fourFunc_wire_382, fourFunc_wire_472});
or_n #(2, 0, 0) OR_95 (fourFunc_wire_231, {fourFunc_wire_384, fourFunc_wire_471});
or_n #(2, 0, 0) OR_96 (fourFunc_wire_227, {fourFunc_wire_386, fourFunc_wire_470});
or_n #(2, 0, 0) OR_97 (fourFunc_wire_223, {fourFunc_wire_388, fourFunc_wire_469});
or_n #(2, 0, 0) OR_98 (fourFunc_wire_219, {fourFunc_wire_390, fourFunc_wire_468});
and_n #(2, 0, 0) AND_195 (fourFunc_wire_210, {fourFunc_wire_507, fourFunc_wire_392_8});
or_n #(2, 0, 0) OR_99 (fourFunc_wire_507, {fourFunc_wire_394, fourFunc_wire_508});
and_n #(2, 0, 0) AND_196 (fourFunc_wire_508, {fourFunc_wire_393, fourFunc_wire_395});
or_n #(2, 0, 0) OR_100 (fourFunc_wire_206, {fourFunc_wire_396, fourFunc_wire_479});
or_n #(2, 0, 0) OR_101 (fourFunc_wire_202, {fourFunc_wire_398, fourFunc_wire_478});
or_n #(2, 0, 0) OR_102 (fourFunc_wire_198, {fourFunc_wire_400, fourFunc_wire_477});
or_n #(2, 0, 0) OR_103 (fourFunc_wire_194, {fourFunc_wire_402, fourFunc_wire_476});
or_n #(2, 0, 0) OR_104 (fourFunc_wire_190, {fourFunc_wire_404, fourFunc_wire_475});
and_n #(2, 0, 0) AND_197 (fourFunc_wire_181, {fourFunc_wire_509, fourFunc_wire_406_8});
or_n #(2, 0, 0) OR_105 (fourFunc_wire_509, {fourFunc_wire_408, fourFunc_wire_510});
and_n #(2, 0, 0) AND_198 (fourFunc_wire_510, {fourFunc_wire_407, fourFunc_wire_409});
or_n #(2, 0, 0) OR_106 (fourFunc_wire_177, {fourFunc_wire_410, fourFunc_wire_486});
or_n #(2, 0, 0) OR_107 (fourFunc_wire_173, {fourFunc_wire_412, fourFunc_wire_485});
or_n #(2, 0, 0) OR_108 (fourFunc_wire_169, {fourFunc_wire_414, fourFunc_wire_484});
or_n #(2, 0, 0) OR_109 (fourFunc_wire_165, {fourFunc_wire_416, fourFunc_wire_483});
or_n #(2, 0, 0) OR_110 (fourFunc_wire_161, {fourFunc_wire_418, fourFunc_wire_482});
and_n #(2, 0, 0) AND_199 (fourFunc_wire_152, {fourFunc_wire_511, fourFunc_wire_420_8});
or_n #(2, 0, 0) OR_111 (fourFunc_wire_511, {fourFunc_wire_422, fourFunc_wire_512});
and_n #(2, 0, 0) AND_200 (fourFunc_wire_512, {fourFunc_wire_421, fourFunc_wire_423});
or_n #(2, 0, 0) OR_112 (fourFunc_wire_147, {fourFunc_wire_424, fourFunc_wire_493});
or_n #(2, 0, 0) OR_113 (fourFunc_wire_142, {fourFunc_wire_426, fourFunc_wire_492});
or_n #(2, 0, 0) OR_114 (fourFunc_wire_137, {fourFunc_wire_428, fourFunc_wire_491});
or_n #(2, 0, 0) OR_115 (fourFunc_wire_132, {fourFunc_wire_430, fourFunc_wire_490});
or_n #(2, 0, 0) OR_116 (fourFunc_wire_127, {fourFunc_wire_432, fourFunc_wire_489});
or_n #(2, 0, 0) OR_117 (fourFunc_wire_93, {fourFunc_wire_513, fourFunc_wire_54_3});
and_n #(2, 0, 0) AND_201 (fourFunc_wire_514, {fourFunc_wire_93_1, fourFunc_wire_515});
notg #(0, 0) NOT_16 (fourFunc_wire_513, fourFunc_wire_53_17);
or_n #(2, 0, 0) OR_118 (fourFunc_wire_88, {fourFunc_wire_516, fourFunc_wire_514});
and_n #(2, 0, 0) AND_202 (fourFunc_wire_517, {fourFunc_wire_88_1, fourFunc_wire_518});
notg #(0, 0) NOT_17 (fourFunc_wire_519, fourFunc_wire_95_25);
or_n #(2, 0, 0) OR_119 (fourFunc_wire_515, {fourFunc_wire_519, fourFunc_wire_94_4});
notg #(0, 0) NOT_18 (fourFunc_wire_520, fourFunc_wire_95_26);
and_n #(2, 0, 0) AND_203 (fourFunc_wire_516, {fourFunc_wire_520, fourFunc_wire_94_5});
or_n #(2, 0, 0) OR_120 (fourFunc_wire_83, {fourFunc_wire_521, fourFunc_wire_517});
and_n #(2, 0, 0) AND_204 (fourFunc_wire_522, {fourFunc_wire_83_1, fourFunc_wire_523});
notg #(0, 0) NOT_19 (fourFunc_wire_524, fourFunc_wire_90_12);
or_n #(2, 0, 0) OR_121 (fourFunc_wire_518, {fourFunc_wire_524, fourFunc_wire_89_4});
notg #(0, 0) NOT_20 (fourFunc_wire_525, fourFunc_wire_90_13);
and_n #(2, 0, 0) AND_205 (fourFunc_wire_521, {fourFunc_wire_525, fourFunc_wire_89_5});
or_n #(2, 0, 0) OR_122 (fourFunc_wire_78, {fourFunc_wire_526, fourFunc_wire_522});
and_n #(2, 0, 0) AND_206 (fourFunc_wire_527, {fourFunc_wire_78_1, fourFunc_wire_528});
notg #(0, 0) NOT_21 (fourFunc_wire_529, fourFunc_wire_85_12);
or_n #(2, 0, 0) OR_123 (fourFunc_wire_523, {fourFunc_wire_529, fourFunc_wire_84_4});
notg #(0, 0) NOT_22 (fourFunc_wire_530, fourFunc_wire_85_13);
and_n #(2, 0, 0) AND_207 (fourFunc_wire_526, {fourFunc_wire_530, fourFunc_wire_84_5});
or_n #(2, 0, 0) OR_124 (fourFunc_wire_73, {fourFunc_wire_531, fourFunc_wire_527});
and_n #(2, 0, 0) AND_208 (fourFunc_wire_532, {fourFunc_wire_73_1, fourFunc_wire_533});
notg #(0, 0) NOT_23 (fourFunc_wire_534, fourFunc_wire_80_12);
or_n #(2, 0, 0) OR_125 (fourFunc_wire_528, {fourFunc_wire_534, fourFunc_wire_79_4});
notg #(0, 0) NOT_24 (fourFunc_wire_535, fourFunc_wire_80_13);
and_n #(2, 0, 0) AND_209 (fourFunc_wire_531, {fourFunc_wire_535, fourFunc_wire_79_5});
or_n #(2, 0, 0) OR_126 (fourFunc_wire_68, {fourFunc_wire_536, fourFunc_wire_532});
and_n #(2, 0, 0) AND_210 (fourFunc_wire_537, {fourFunc_wire_68_1, fourFunc_wire_538});
notg #(0, 0) NOT_25 (fourFunc_wire_539, fourFunc_wire_75_12);
or_n #(2, 0, 0) OR_127 (fourFunc_wire_533, {fourFunc_wire_539, fourFunc_wire_74_4});
notg #(0, 0) NOT_26 (fourFunc_wire_540, fourFunc_wire_75_13);
and_n #(2, 0, 0) AND_211 (fourFunc_wire_536, {fourFunc_wire_540, fourFunc_wire_74_5});
or_n #(2, 0, 0) OR_128 (fourFunc_wire_63, {fourFunc_wire_541, fourFunc_wire_537});
and_n #(2, 0, 0) AND_212 (fourFunc_wire_542, {fourFunc_wire_63_1, fourFunc_wire_543});
notg #(0, 0) NOT_27 (fourFunc_wire_544, fourFunc_wire_70_12);
or_n #(2, 0, 0) OR_129 (fourFunc_wire_538, {fourFunc_wire_544, fourFunc_wire_69_4});
notg #(0, 0) NOT_28 (fourFunc_wire_545, fourFunc_wire_70_13);
and_n #(2, 0, 0) AND_213 (fourFunc_wire_541, {fourFunc_wire_545, fourFunc_wire_69_5});
or_n #(2, 0, 0) OR_130 (fourFunc_wire_57, {fourFunc_wire_60_1, fourFunc_wire_59_3});
or_n #(2, 0, 0) OR_131 (fourFunc_wire_60, {fourFunc_wire_546, fourFunc_wire_542});
notg #(0, 0) NOT_29 (fourFunc_wire_547, fourFunc_wire_65_12);
or_n #(2, 0, 0) OR_132 (fourFunc_wire_543, {fourFunc_wire_547, fourFunc_wire_64_4});
notg #(0, 0) NOT_30 (fourFunc_wire_548, fourFunc_wire_65_13);
and_n #(2, 0, 0) AND_214 (fourFunc_wire_546, {fourFunc_wire_548, fourFunc_wire_64_5});
bufg #(0, 0) BUF_1 (fourFunc_wire_549, 1'b0);
and_n #(2, 0, 0) AND_215 (fourFunc_wire_560, {fourFunc_wire_96, fourFunc_wire_551_0});
and_n #(2, 0, 0) AND_216 (fourFunc_wire_561, {fourFunc_wire_119, fourFunc_wire_551_1});
and_n #(2, 0, 0) AND_217 (fourFunc_wire_562, {fourFunc_wire_116, fourFunc_wire_551_2});
and_n #(2, 0, 0) AND_218 (fourFunc_wire_563, {fourFunc_wire_113, fourFunc_wire_551_3});
and_n #(2, 0, 0) AND_219 (fourFunc_wire_564, {fourFunc_wire_110, fourFunc_wire_551_4});
and_n #(2, 0, 0) AND_220 (fourFunc_wire_565, {fourFunc_wire_107, fourFunc_wire_551_5});
and_n #(2, 0, 0) AND_221 (fourFunc_wire_566, {fourFunc_wire_104, fourFunc_wire_551_6});
and_n #(2, 0, 0) AND_222 (fourFunc_wire_567, {fourFunc_wire_101, fourFunc_wire_551_7});
and_n #(2, 0, 0) AND_223 (fourFunc_wire_568, {fourFunc_wire_97, fourFunc_wire_551_8});
and_n #(2, 0, 0) AND_224 (fourFunc_wire_569, {fourFunc_wire_99, fourFunc_wire_551_9});
notg #(0, 0) NOT_31 (fourFunc_wire_570, fourFunc_wire_551_10);
notg #(0, 0) NOT_32 (fourFunc_wire_571, fourFunc_wire_551_11);
notg #(0, 0) NOT_33 (fourFunc_wire_572, fourFunc_wire_551_12);
notg #(0, 0) NOT_34 (fourFunc_wire_573, fourFunc_wire_551_13);
notg #(0, 0) NOT_35 (fourFunc_wire_574, fourFunc_wire_551_14);
notg #(0, 0) NOT_36 (fourFunc_wire_575, fourFunc_wire_551_15);
notg #(0, 0) NOT_37 (fourFunc_wire_576, fourFunc_wire_551_16);
notg #(0, 0) NOT_38 (fourFunc_wire_577, fourFunc_wire_551_17);
notg #(0, 0) NOT_39 (fourFunc_wire_578, fourFunc_wire_551_18);
notg #(0, 0) NOT_40 (fourFunc_wire_579, fourFunc_wire_551_19);
or_n #(2, 0, 0) OR_133 (fourFunc_wire_580, {fourFunc_wire_570, fourFunc_wire_581_0});
or_n #(2, 0, 0) OR_134 (fourFunc_wire_582, {fourFunc_wire_583, fourFunc_wire_581_1});
notg #(0, 0) NOT_41 (fourFunc_wire_584, fourFunc_wire_585);
and_n #(2, 0, 0) AND_225 (fourFunc_wire_583, {fourFunc_wire_584, fourFunc_wire_586_0});
or_n #(4, 0, 0) OR_135 (fourFunc_wire_587, {fourFunc_wire_588_0, fourFunc_wire_589_0, fourFunc_wire_590_0, fourFunc_wire_586_1});
and_n #(2, 0, 0) AND_226 (fourFunc_wire_50, {fourFunc_wire_2_8, fourFunc_wire_8_10});
notg #(0, 0) NOT_42 (fourFunc_wire_600, fourFunc_wire_2_9);
and_n #(2, 0, 0) AND_227 (fourFunc_wire_601, {fourFunc_wire_602, fourFunc_wire_603});
or_n #(2, 0, 0) OR_136 (fourFunc_wire_603, {fourFunc_wire_600, fourFunc_wire_604_0});
notg #(0, 0) NOT_43 (fourFunc_wire_602, fourFunc_wire_599_0);
or_n #(3, 0, 0) OR_137 (fourFunc_wire_605, {fourFunc_wire_604_1, fourFunc_wire_589_1, fourFunc_wire_599_1});
and_n #(2, 0, 0) AND_228 (fourFunc_wire_606, {fourFunc_wire_607, fourFunc_wire_51});
notg #(0, 0) NOT_44 (fourFunc_wire_607, fourFunc_wire_608_0);
or_n #(2, 0, 0) OR_138 (fourFunc_wire_609, {fourFunc_wire_608_1, fourFunc_wire_589_2});
and_n #(2, 0, 0) AND_229 (fourFunc_wire_48, {fourFunc_wire_3_7, fourFunc_wire_50_1});
and_n #(2, 0, 0) AND_230 (fourFunc_wire_610, {fourFunc_wire_611, fourFunc_wire_49});
notg #(0, 0) NOT_45 (fourFunc_wire_611, fourFunc_wire_608_2);
and_n #(2, 0, 0) AND_231 (fourFunc_wire_612, {fourFunc_wire_10_8, fourFunc_wire_588_1});
notg #(0, 0) NOT_46 (fourFunc_wire_613, fourFunc_wire_10_9);
and_n #(2, 0, 0) AND_232 (fourFunc_wire_614, {fourFunc_wire_615, fourFunc_wire_47});
notg #(0, 0) NOT_47 (fourFunc_wire_615, fourFunc_wire_608_3);
or_n #(2, 0, 0) OR_139 (fourFunc_wire_608, {fourFunc_wire_604_2, fourFunc_wire_599_2});
notg #(0, 0) NOT_48 (fourFunc_wire_616, fourFunc_wire_9_7);
and_n #(2, 0, 0) AND_233 (fourFunc_wire_617, {fourFunc_wire_9_8, fourFunc_wire_604_3});
notg #(0, 0) NOT_49 (fourFunc_wire_618, fourFunc_wire_9_9);
notg #(0, 0) NOT_50 (fourFunc_wire_619, fourFunc_wire_9_10);
notg #(0, 0) NOT_51 (fourFunc_wire_620, fourFunc_wire_9_11);
notg #(0, 0) NOT_52 (fourFunc_wire_621, fourFunc_wire_9_12);
notg #(0, 0) NOT_53 (fourFunc_wire_622, fourFunc_wire_9_13);
notg #(0, 0) NOT_54 (fourFunc_wire_623, fourFunc_wire_9_14);
notg #(0, 0) NOT_55 (fourFunc_wire_624, fourFunc_wire_9_15);
or_n #(2, 0, 0) OR_140 (fourFunc_wire_625, {fourFunc_wire_9_16, fourFunc_wire_626_0});
or_n #(2, 0, 0) OR_141 (fourFunc_wire_627, {fourFunc_wire_9_17, fourFunc_wire_628_0});
or_n #(2, 0, 0) OR_142 (fourFunc_wire_629, {fourFunc_wire_9_18, fourFunc_wire_630_0});
or_n #(2, 0, 0) OR_143 (fourFunc_wire_631, {fourFunc_wire_9_19, fourFunc_wire_632_0});
or_n #(2, 0, 0) OR_144 (fourFunc_wire_633, {fourFunc_wire_9_20, fourFunc_wire_634_0});
or_n #(2, 0, 0) OR_145 (fourFunc_wire_635, {fourFunc_wire_9_21, fourFunc_wire_636_0});
or_n #(2, 0, 0) OR_146 (fourFunc_wire_637, {fourFunc_wire_9_22, fourFunc_wire_638_0});
or_n #(2, 0, 0) OR_147 (fourFunc_wire_639, {fourFunc_wire_9_23, fourFunc_wire_640_0});
and_n #(2, 0, 0) AND_234 (fourFunc_wire_604, {fourFunc_wire_581_2, fourFunc_wire_641_0});
notg #(0, 0) NOT_56 (fourFunc_wire_642, fourFunc_wire_604_4);
and_n #(2, 0, 0) AND_235 (fourFunc_wire_643, {fourFunc_wire_604_5, fourFunc_wire_628_1});
notg #(0, 0) NOT_57 (fourFunc_wire_644, fourFunc_wire_604_6);
notg #(0, 0) NOT_58 (fourFunc_wire_645, fourFunc_wire_604_7);
notg #(0, 0) NOT_59 (fourFunc_wire_646, fourFunc_wire_604_8);
and_n #(2, 0, 0) AND_236 (fourFunc_wire_647, {fourFunc_wire_604_9, fourFunc_wire_626_1});
or_n #(3, 0, 0) OR_148 (fourFunc_wire_648, {fourFunc_wire_604_10, fourFunc_wire_588_2, fourFunc_wire_599_3});
notg #(0, 0) NOT_60 (fourFunc_wire_649, fourFunc_wire_604_11);
and_n #(2, 0, 0) AND_237 (fourFunc_wire_650, {fourFunc_wire_604_12, fourFunc_wire_634_1});
notg #(0, 0) NOT_61 (fourFunc_wire_651, fourFunc_wire_604_13);
and_n #(2, 0, 0) AND_238 (fourFunc_wire_652, {fourFunc_wire_604_14, fourFunc_wire_636_1});
notg #(0, 0) NOT_62 (fourFunc_wire_653, fourFunc_wire_604_15);
and_n #(2, 0, 0) AND_239 (fourFunc_wire_654, {fourFunc_wire_604_16, fourFunc_wire_630_1});
notg #(0, 0) NOT_63 (fourFunc_wire_655, fourFunc_wire_604_17);
and_n #(2, 0, 0) AND_240 (fourFunc_wire_656, {fourFunc_wire_604_18, fourFunc_wire_640_1});
notg #(0, 0) NOT_64 (fourFunc_wire_657, fourFunc_wire_604_19);
and_n #(2, 0, 0) AND_241 (fourFunc_wire_658, {fourFunc_wire_604_20, fourFunc_wire_632_1});
notg #(0, 0) NOT_65 (fourFunc_wire_659, fourFunc_wire_604_21);
and_n #(2, 0, 0) AND_242 (fourFunc_wire_660, {fourFunc_wire_604_22, fourFunc_wire_638_1});
notg #(0, 0) NOT_66 (fourFunc_wire_661, fourFunc_wire_604_23);
and_n #(2, 0, 0) AND_243 (fourFunc_wire_662, {fourFunc_wire_604_24, fourFunc_wire_625});
notg #(0, 0) NOT_67 (fourFunc_wire_663, fourFunc_wire_604_25);
and_n #(2, 0, 0) AND_244 (fourFunc_wire_664, {fourFunc_wire_604_26, fourFunc_wire_627});
notg #(0, 0) NOT_68 (fourFunc_wire_665, fourFunc_wire_604_27);
and_n #(2, 0, 0) AND_245 (fourFunc_wire_666, {fourFunc_wire_604_28, fourFunc_wire_629});
notg #(0, 0) NOT_69 (fourFunc_wire_667, fourFunc_wire_604_29);
and_n #(2, 0, 0) AND_246 (fourFunc_wire_668, {fourFunc_wire_604_30, fourFunc_wire_631});
notg #(0, 0) NOT_70 (fourFunc_wire_669, fourFunc_wire_604_31);
and_n #(2, 0, 0) AND_247 (fourFunc_wire_670, {fourFunc_wire_604_32, fourFunc_wire_633});
notg #(0, 0) NOT_71 (fourFunc_wire_671, fourFunc_wire_604_33);
and_n #(2, 0, 0) AND_248 (fourFunc_wire_672, {fourFunc_wire_604_34, fourFunc_wire_635});
notg #(0, 0) NOT_72 (fourFunc_wire_673, fourFunc_wire_604_35);
and_n #(2, 0, 0) AND_249 (fourFunc_wire_674, {fourFunc_wire_604_36, fourFunc_wire_637});
notg #(0, 0) NOT_73 (fourFunc_wire_675, fourFunc_wire_604_37);
and_n #(2, 0, 0) AND_250 (fourFunc_wire_676, {fourFunc_wire_604_38, fourFunc_wire_639});
or_n #(2, 0, 0) OR_149 (fourFunc_wire_434, {fourFunc_wire_677, fourFunc_wire_678});
and_n #(2, 0, 0) AND_251 (fourFunc_wire_677, {fourFunc_wire_586_2, fourFunc_wire_40});
notg #(0, 0) NOT_74 (fourFunc_wire_679, fourFunc_wire_586_3);
and_n #(2, 0, 0) AND_252 (fourFunc_wire_678, {fourFunc_wire_679, fourFunc_wire_552_0});
or_n #(2, 0, 0) OR_150 (fourFunc_wire_446, {fourFunc_wire_680, fourFunc_wire_681});
and_n #(2, 0, 0) AND_253 (fourFunc_wire_680, {fourFunc_wire_586_4, fourFunc_wire_4});
notg #(0, 0) NOT_75 (fourFunc_wire_682, fourFunc_wire_586_5);
and_n #(2, 0, 0) AND_254 (fourFunc_wire_681, {fourFunc_wire_682, fourFunc_wire_553_0});
or_n #(2, 0, 0) OR_151 (fourFunc_wire_350, {fourFunc_wire_683, fourFunc_wire_684});
and_n #(2, 0, 0) AND_255 (fourFunc_wire_683, {fourFunc_wire_586_6, fourFunc_wire_42});
notg #(0, 0) NOT_76 (fourFunc_wire_685, fourFunc_wire_586_7);
and_n #(2, 0, 0) AND_256 (fourFunc_wire_684, {fourFunc_wire_685, fourFunc_wire_554_0});
or_n #(2, 0, 0) OR_152 (fourFunc_wire_364, {fourFunc_wire_686, fourFunc_wire_687});
and_n #(2, 0, 0) AND_257 (fourFunc_wire_686, {fourFunc_wire_586_8, fourFunc_wire_12});
notg #(0, 0) NOT_77 (fourFunc_wire_688, fourFunc_wire_586_9);
and_n #(2, 0, 0) AND_258 (fourFunc_wire_687, {fourFunc_wire_688, fourFunc_wire_555_0});
or_n #(2, 0, 0) OR_153 (fourFunc_wire_378, {fourFunc_wire_689, fourFunc_wire_690});
and_n #(2, 0, 0) AND_259 (fourFunc_wire_689, {fourFunc_wire_586_10, fourFunc_wire_25});
notg #(0, 0) NOT_78 (fourFunc_wire_691, fourFunc_wire_586_11);
and_n #(2, 0, 0) AND_260 (fourFunc_wire_690, {fourFunc_wire_691, fourFunc_wire_556_0});
and_n #(2, 0, 0) AND_261 (fourFunc_wire_392, {fourFunc_wire_692, fourFunc_wire_557_0});
notg #(0, 0) NOT_79 (fourFunc_wire_692, fourFunc_wire_586_12);
and_n #(2, 0, 0) AND_262 (fourFunc_wire_406, {fourFunc_wire_693, fourFunc_wire_558_0});
notg #(0, 0) NOT_80 (fourFunc_wire_693, fourFunc_wire_586_13);
or_n #(2, 0, 0) OR_154 (fourFunc_wire_420, {fourFunc_wire_694, fourFunc_wire_695});
and_n #(2, 0, 0) AND_263 (fourFunc_wire_694, {fourFunc_wire_586_14, fourFunc_wire_17});
notg #(0, 0) NOT_81 (fourFunc_wire_696, fourFunc_wire_586_15);
and_n #(2, 0, 0) AND_264 (fourFunc_wire_695, {fourFunc_wire_696, fourFunc_wire_559_0});
and_n #(2, 0, 0) AND_265 (fourFunc_wire_697, {fourFunc_wire_145, fourFunc_wire_665});
and_n #(2, 0, 0) AND_266 (fourFunc_wire_698, {fourFunc_wire_140, fourFunc_wire_669});
and_n #(2, 0, 0) AND_267 (fourFunc_wire_699, {fourFunc_wire_135, fourFunc_wire_671});
and_n #(2, 0, 0) AND_268 (fourFunc_wire_700, {fourFunc_wire_130, fourFunc_wire_667});
and_n #(2, 0, 0) AND_269 (fourFunc_wire_701, {fourFunc_wire_125, fourFunc_wire_673});
and_n #(2, 0, 0) AND_270 (fourFunc_wire_702, {fourFunc_wire_155, fourFunc_wire_661});
and_n #(2, 0, 0) AND_271 (fourFunc_wire_703, {fourFunc_wire_150, fourFunc_wire_663});
or_n #(2, 0, 0) OR_155 (fourFunc_wire_704, {fourFunc_wire_592, fourFunc_wire_599_4});
and_n #(2, 0, 0) AND_272 (fourFunc_wire_591, {fourFunc_wire_612, fourFunc_wire_705});
notg #(0, 0) NOT_82 (fourFunc_wire_705, fourFunc_wire_598_0);
and_n #(2, 0, 0) AND_273 (fourFunc_wire_706, {fourFunc_wire_588_3, fourFunc_wire_613});
notg #(0, 0) NOT_83 (fourFunc_wire_707, fourFunc_wire_598_1);
and_n #(2, 0, 0) AND_274 (fourFunc_wire_593, {fourFunc_wire_707, fourFunc_wire_589_3});
notg #(0, 0) NOT_84 (fourFunc_wire_708, fourFunc_wire_598_2);
and_n #(2, 0, 0) AND_275 (fourFunc_wire_594, {fourFunc_wire_708, fourFunc_wire_590_1});
notg #(0, 0) NOT_85 (fourFunc_wire_709, fourFunc_wire_598_3);
and_n #(2, 0, 0) AND_276 (fourFunc_wire_595, {fourFunc_wire_709, fourFunc_wire_586_16});
and_n #(2, 0, 0) AND_277 (fourFunc_wire_710, {fourFunc_wire_581_3, fourFunc_wire_641_1});
or_n #(2, 0, 0) OR_156 (fourFunc_wire_711, {fourFunc_wire_710, fourFunc_wire_706});
notg #(0, 0) NOT_86 (fourFunc_wire_712, fourFunc_wire_598_4);
and_n #(2, 0, 0) AND_278 (fourFunc_wire_596, {fourFunc_wire_712, fourFunc_wire_711});
and_n #(2, 0, 0) AND_279 (fourFunc_wire_713, {fourFunc_wire_581_4, fourFunc_wire_714});
or_n #(2, 0, 0) OR_157 (fourFunc_wire_715, {fourFunc_wire_704, fourFunc_wire_713});
notg #(0, 0) NOT_87 (fourFunc_wire_714, fourFunc_wire_641_2);
notg #(0, 0) NOT_88 (fourFunc_wire_716, fourFunc_wire_598_5);
and_n #(2, 0, 0) AND_280 (fourFunc_wire_597, {fourFunc_wire_716, fourFunc_wire_715});
or_n #(2, 0, 0) OR_158 (fourFunc_wire_717, {fourFunc_wire_599_5, fourFunc_wire_718});
notg #(0, 0) NOT_89 (fourFunc_wire_719, fourFunc_wire_599_6);
notg #(0, 0) NOT_90 (fourFunc_wire_720, fourFunc_wire_599_7);
notg #(0, 0) NOT_91 (fourFunc_wire_721, fourFunc_wire_599_8);
notg #(0, 0) NOT_92 (fourFunc_wire_722, fourFunc_wire_599_9);
notg #(0, 0) NOT_93 (fourFunc_wire_723, fourFunc_wire_599_10);
notg #(0, 0) NOT_94 (fourFunc_wire_724, fourFunc_wire_599_11);
notg #(0, 0) NOT_95 (fourFunc_wire_725, fourFunc_wire_599_12);
notg #(0, 0) NOT_96 (fourFunc_wire_726, fourFunc_wire_599_13);
notg #(0, 0) NOT_97 (fourFunc_wire_727, fourFunc_wire_599_14);
notg #(0, 0) NOT_98 (fourFunc_wire_728, fourFunc_wire_599_15);
notg #(0, 0) NOT_99 (fourFunc_wire_729, fourFunc_wire_599_16);
notg #(0, 0) NOT_100 (fourFunc_wire_730, fourFunc_wire_599_17);
notg #(0, 0) NOT_101 (fourFunc_wire_731, fourFunc_wire_599_18);
notg #(0, 0) NOT_102 (fourFunc_wire_732, fourFunc_wire_599_19);
notg #(0, 0) NOT_103 (fourFunc_wire_733, fourFunc_wire_599_20);
notg #(0, 0) NOT_104 (fourFunc_wire_734, fourFunc_wire_599_21);
notg #(0, 0) NOT_105 (fourFunc_wire_735, fourFunc_wire_599_22);
notg #(0, 0) NOT_106 (fourFunc_wire_736, fourFunc_wire_599_23);
notg #(0, 0) NOT_107 (fourFunc_wire_737, fourFunc_wire_599_24);
notg #(0, 0) NOT_108 (fourFunc_wire_738, fourFunc_wire_599_25);
notg #(0, 0) NOT_109 (fourFunc_wire_739, fourFunc_wire_599_26);
notg #(0, 0) NOT_110 (fourFunc_wire_740, fourFunc_wire_599_27);
notg #(0, 0) NOT_111 (fourFunc_wire_741, fourFunc_wire_599_28);
notg #(0, 0) NOT_112 (fourFunc_wire_742, fourFunc_wire_599_29);
notg #(0, 0) NOT_113 (fourFunc_wire_743, fourFunc_wire_599_30);
notg #(0, 0) NOT_114 (fourFunc_wire_744, fourFunc_wire_599_31);
and_n #(2, 0, 0) AND_281 (fourFunc_wire_745, {fourFunc_wire_719, fourFunc_wire_626_2});
and_n #(2, 0, 0) AND_282 (fourFunc_wire_746, {fourFunc_wire_720, fourFunc_wire_628_2});
and_n #(2, 0, 0) AND_283 (fourFunc_wire_747, {fourFunc_wire_721, fourFunc_wire_630_2});
and_n #(2, 0, 0) AND_284 (fourFunc_wire_748, {fourFunc_wire_722, fourFunc_wire_634_2});
and_n #(2, 0, 0) AND_285 (fourFunc_wire_749, {fourFunc_wire_723, fourFunc_wire_636_2});
and_n #(2, 0, 0) AND_286 (fourFunc_wire_750, {fourFunc_wire_724, fourFunc_wire_632_2});
and_n #(2, 0, 0) AND_287 (fourFunc_wire_751, {fourFunc_wire_725, fourFunc_wire_638_2});
and_n #(2, 0, 0) AND_288 (fourFunc_wire_752, {fourFunc_wire_726, fourFunc_wire_640_2});
and_n #(2, 0, 0) AND_289 (fourFunc_wire_753, {fourFunc_wire_754, fourFunc_wire_730});
or_n #(2, 0, 0) OR_159 (fourFunc_wire_755, {fourFunc_wire_560, fourFunc_wire_756});
and_n #(2, 0, 0) AND_290 (fourFunc_wire_757, {fourFunc_wire_755, fourFunc_wire_646});
or_n #(2, 0, 0) OR_160 (fourFunc_wire_754, {fourFunc_wire_757, fourFunc_wire_758});
nor_n #(2, 0, 0) NOR_3 (fourFunc_wire_756, {fourFunc_wire_551_20, fourFunc_wire_52});
and_n #(2, 0, 0) AND_291 (fourFunc_wire_758, {fourFunc_wire_647, fourFunc_wire_618});
and_n #(2, 0, 0) AND_292 (fourFunc_wire_759, {fourFunc_wire_760, fourFunc_wire_727});
or_n #(2, 0, 0) OR_161 (fourFunc_wire_761, {fourFunc_wire_561, fourFunc_wire_762});
and_n #(2, 0, 0) AND_293 (fourFunc_wire_763, {fourFunc_wire_642, fourFunc_wire_761});
or_n #(2, 0, 0) OR_162 (fourFunc_wire_760, {fourFunc_wire_763, fourFunc_wire_764});
and_n #(2, 0, 0) AND_294 (fourFunc_wire_762, {fourFunc_wire_571, fourFunc_wire_91});
and_n #(2, 0, 0) AND_295 (fourFunc_wire_764, {fourFunc_wire_643, fourFunc_wire_616});
and_n #(2, 0, 0) AND_296 (fourFunc_wire_765, {fourFunc_wire_766, fourFunc_wire_733});
or_n #(2, 0, 0) OR_163 (fourFunc_wire_767, {fourFunc_wire_562, fourFunc_wire_768});
and_n #(2, 0, 0) AND_297 (fourFunc_wire_769, {fourFunc_wire_653, fourFunc_wire_767});
or_n #(2, 0, 0) OR_164 (fourFunc_wire_766, {fourFunc_wire_769, fourFunc_wire_770});
and_n #(2, 0, 0) AND_298 (fourFunc_wire_768, {fourFunc_wire_576, fourFunc_wire_86});
and_n #(2, 0, 0) AND_299 (fourFunc_wire_770, {fourFunc_wire_654, fourFunc_wire_621});
and_n #(2, 0, 0) AND_300 (fourFunc_wire_771, {fourFunc_wire_772, fourFunc_wire_731});
or_n #(2, 0, 0) OR_165 (fourFunc_wire_773, {fourFunc_wire_563, fourFunc_wire_774});
and_n #(2, 0, 0) AND_301 (fourFunc_wire_775, {fourFunc_wire_649, fourFunc_wire_773});
or_n #(2, 0, 0) OR_166 (fourFunc_wire_772, {fourFunc_wire_775, fourFunc_wire_776});
and_n #(2, 0, 0) AND_302 (fourFunc_wire_774, {fourFunc_wire_574, fourFunc_wire_81});
and_n #(2, 0, 0) AND_303 (fourFunc_wire_776, {fourFunc_wire_650, fourFunc_wire_619});
and_n #(2, 0, 0) AND_304 (fourFunc_wire_777, {fourFunc_wire_778, fourFunc_wire_732});
or_n #(2, 0, 0) OR_167 (fourFunc_wire_779, {fourFunc_wire_564, fourFunc_wire_780});
and_n #(2, 0, 0) AND_305 (fourFunc_wire_781, {fourFunc_wire_651, fourFunc_wire_779});
or_n #(2, 0, 0) OR_168 (fourFunc_wire_778, {fourFunc_wire_781, fourFunc_wire_782});
and_n #(2, 0, 0) AND_306 (fourFunc_wire_780, {fourFunc_wire_575, fourFunc_wire_76});
and_n #(2, 0, 0) AND_307 (fourFunc_wire_782, {fourFunc_wire_652, fourFunc_wire_620});
and_n #(2, 0, 0) AND_308 (fourFunc_wire_783, {fourFunc_wire_784, fourFunc_wire_735});
or_n #(2, 0, 0) OR_169 (fourFunc_wire_785, {fourFunc_wire_565, fourFunc_wire_786});
and_n #(2, 0, 0) AND_309 (fourFunc_wire_787, {fourFunc_wire_657, fourFunc_wire_785});
or_n #(2, 0, 0) OR_170 (fourFunc_wire_784, {fourFunc_wire_787, fourFunc_wire_788});
and_n #(2, 0, 0) AND_310 (fourFunc_wire_786, {fourFunc_wire_578, fourFunc_wire_71});
and_n #(2, 0, 0) AND_311 (fourFunc_wire_788, {fourFunc_wire_658, fourFunc_wire_623});
and_n #(2, 0, 0) AND_312 (fourFunc_wire_789, {fourFunc_wire_790, fourFunc_wire_736});
or_n #(2, 0, 0) OR_171 (fourFunc_wire_791, {fourFunc_wire_566, fourFunc_wire_792});
and_n #(2, 0, 0) AND_313 (fourFunc_wire_793, {fourFunc_wire_659, fourFunc_wire_791});
or_n #(2, 0, 0) OR_172 (fourFunc_wire_790, {fourFunc_wire_793, fourFunc_wire_794});
and_n #(2, 0, 0) AND_314 (fourFunc_wire_792, {fourFunc_wire_579, fourFunc_wire_66});
and_n #(2, 0, 0) AND_315 (fourFunc_wire_794, {fourFunc_wire_660, fourFunc_wire_624});
and_n #(2, 0, 0) AND_316 (fourFunc_wire_795, {fourFunc_wire_796, fourFunc_wire_734});
or_n #(2, 0, 0) OR_173 (fourFunc_wire_797, {fourFunc_wire_567, fourFunc_wire_798});
and_n #(2, 0, 0) AND_317 (fourFunc_wire_799, {fourFunc_wire_655, fourFunc_wire_797});
or_n #(2, 0, 0) OR_174 (fourFunc_wire_796, {fourFunc_wire_799, fourFunc_wire_800});
and_n #(2, 0, 0) AND_318 (fourFunc_wire_798, {fourFunc_wire_577, fourFunc_wire_61});
and_n #(2, 0, 0) AND_319 (fourFunc_wire_800, {fourFunc_wire_656, fourFunc_wire_622});
and_n #(2, 0, 0) AND_320 (fourFunc_wire_801, {fourFunc_wire_728, fourFunc_wire_802});
or_n #(2, 0, 0) OR_175 (fourFunc_wire_802, {fourFunc_wire_617, fourFunc_wire_803});
or_n #(2, 0, 0) OR_176 (fourFunc_wire_804, {fourFunc_wire_568, fourFunc_wire_805});
and_n #(2, 0, 0) AND_321 (fourFunc_wire_805, {fourFunc_wire_572, fourFunc_wire_58});
and_n #(2, 0, 0) AND_322 (fourFunc_wire_803, {fourFunc_wire_644, fourFunc_wire_804});
and_n #(3, 0, 0) AND_323 (fourFunc_wire_806, {fourFunc_wire_729, fourFunc_wire_645, fourFunc_wire_807});
or_n #(2, 0, 0) OR_177 (fourFunc_wire_807, {fourFunc_wire_569, fourFunc_wire_808});
and_n #(2, 0, 0) AND_324 (fourFunc_wire_808, {fourFunc_wire_573, fourFunc_wire_55});
and_n #(2, 0, 0) AND_325 (fourFunc_wire_809, {fourFunc_wire_737, fourFunc_wire_810});
or_n #(2, 0, 0) OR_178 (fourFunc_wire_810, {fourFunc_wire_662, fourFunc_wire_702});
notg #(0, 0) NOT_115 (fourFunc_wire_718, fourFunc_wire_811);
and_n #(2, 0, 0) AND_326 (fourFunc_wire_812, {fourFunc_wire_738, fourFunc_wire_813});
or_n #(2, 0, 0) OR_179 (fourFunc_wire_813, {fourFunc_wire_664, fourFunc_wire_703});
and_n #(2, 0, 0) AND_327 (fourFunc_wire_814, {fourFunc_wire_739, fourFunc_wire_815});
or_n #(2, 0, 0) OR_180 (fourFunc_wire_815, {fourFunc_wire_666, fourFunc_wire_697});
and_n #(2, 0, 0) AND_328 (fourFunc_wire_816, {fourFunc_wire_741, fourFunc_wire_817});
or_n #(2, 0, 0) OR_181 (fourFunc_wire_817, {fourFunc_wire_670, fourFunc_wire_698});
and_n #(2, 0, 0) AND_329 (fourFunc_wire_818, {fourFunc_wire_742, fourFunc_wire_819});
or_n #(2, 0, 0) OR_182 (fourFunc_wire_819, {fourFunc_wire_672, fourFunc_wire_699});
and_n #(2, 0, 0) AND_330 (fourFunc_wire_820, {fourFunc_wire_740, fourFunc_wire_821});
or_n #(2, 0, 0) OR_183 (fourFunc_wire_821, {fourFunc_wire_668, fourFunc_wire_700});
and_n #(2, 0, 0) AND_331 (fourFunc_wire_822, {fourFunc_wire_743, fourFunc_wire_823});
or_n #(2, 0, 0) OR_184 (fourFunc_wire_823, {fourFunc_wire_674, fourFunc_wire_701});
and_n #(2, 0, 0) AND_332 (fourFunc_wire_824, {fourFunc_wire_825, fourFunc_wire_744});
or_n #(2, 0, 0) OR_185 (fourFunc_wire_825, {fourFunc_wire_676, fourFunc_wire_826});
or_n #(2, 0, 0) OR_186 (fourFunc_wire_827, {fourFunc_wire_499, fourFunc_wire_487});
and_n #(2, 0, 0) AND_333 (fourFunc_wire_826, {fourFunc_wire_675, fourFunc_wire_827});
nor_n #(4, 0, 0) NOR_4 (fourFunc_wire_811, {fourFunc_wire_604_39, fourFunc_wire_590_2, fourFunc_wire_589_4, fourFunc_wire_586_17});
bufg #(0, 0) BUF_2 (busy_net_0, fourFunc_wire_587);
bufg #(0, 0) BUF_3 (fourFunc_wire_550, clk_net_0);
bufg #(0, 0) BUF_4 (fourFunc_wire_9, func_1);
bufg #(0, 0) BUF_5 (fourFunc_wire_585, func_0);
bufg #(0, 0) BUF_6 (resultFPart_7, fourFunc_wire_54_4);
bufg #(0, 0) BUF_7 (resultFPart_6, fourFunc_wire_94_6);
bufg #(0, 0) BUF_8 (resultFPart_5, fourFunc_wire_89_6);
bufg #(0, 0) BUF_9 (resultFPart_4, fourFunc_wire_84_6);
bufg #(0, 0) BUF_10 (resultFPart_3, fourFunc_wire_79_6);
bufg #(0, 0) BUF_11 (resultFPart_2, fourFunc_wire_74_6);
bufg #(0, 0) BUF_12 (resultFPart_1, fourFunc_wire_69_6);
bufg #(0, 0) BUF_13 (resultFPart_0, fourFunc_wire_64_6);
bufg #(0, 0) BUF_14 (resultIPart_1, fourFunc_wire_59_4);
bufg #(0, 0) BUF_15 (resultIPart_0, fourFunc_wire_56_2);
bufg #(0, 0) BUF_16 (fourFunc_wire_598, rst_net_0);
bufg #(0, 0) BUF_17 (fourFunc_wire_641, start_net_0);
bufg #(0, 0) BUF_18 (fourFunc_wire_626, x_7);
bufg #(0, 0) BUF_19 (fourFunc_wire_628, x_6);
bufg #(0, 0) BUF_20 (fourFunc_wire_630, x_5);
bufg #(0, 0) BUF_21 (fourFunc_wire_634, x_4);
bufg #(0, 0) BUF_22 (fourFunc_wire_636, x_3);
bufg #(0, 0) BUF_23 (fourFunc_wire_632, x_2);
bufg #(0, 0) BUF_24 (fourFunc_wire_638, x_1);
bufg #(0, 0) BUF_25 (fourFunc_wire_640, x_0);
and_n #(2, 0, 0) AND_334 (NOT_intermediateXXXwire_676_AND_intermediateXXXwire_673, {fourFunc_wire_551_21, NOT_intermediateXXXwire_676});
and_n #(2, 0, 0) AND_335 (fourFunc_wire_828, {fourFunc_wire_582_0, fourFunc_wire_580});
or_n #(2, 0, 0) OR_187 (NOT_intermediateXXXwire_676_AND_intermediateXXXwire_673_OR_intermediateXXXwire_676_AND_intermediateXXXwire_674, {NOT_intermediateXXXwire_676_AND_intermediateXXXwire_673, fourFunc_wire_828});
notg #(0, 0) NOT_116 (NOT_intermediateXXXwire_676, fourFunc_wire_582_1);
and_n #(2, 0, 0) AND_336 (NOT_intermediateXXXwire_686_AND_intermediateXXXwire_14, {fourFunc_wire_2_10, NOT_intermediateXXXwire_686});
and_n #(2, 0, 0) AND_337 (fourFunc_wire_829, {fourFunc_wire_605_0, fourFunc_wire_601});
or_n #(2, 0, 0) OR_188 (NOT_intermediateXXXwire_686_AND_intermediateXXXwire_14_OR_intermediateXXXwire_686_AND_intermediateXXXwire_682, {NOT_intermediateXXXwire_686_AND_intermediateXXXwire_14, fourFunc_wire_829});
notg #(0, 0) NOT_117 (NOT_intermediateXXXwire_686, fourFunc_wire_605_1);
and_n #(2, 0, 0) AND_338 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_17, {fourFunc_wire_10_10, NOT_intermediateXXXwire_690_0});
and_n #(2, 0, 0) AND_339 (fourFunc_wire_830, {fourFunc_wire_609_0, fourFunc_wire_614});
or_n #(2, 0, 0) OR_189 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_17_OR_intermediateXXXwire_690_AND_intermediateXXXwire_695, {NOT_intermediateXXXwire_690_AND_intermediateXXXwire_17, fourFunc_wire_830});
notg #(0, 0) NOT_118 (NOT_intermediateXXXwire_690, fourFunc_wire_609_1);
and_n #(2, 0, 0) AND_340 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_16, {fourFunc_wire_3_8, NOT_intermediateXXXwire_690_1});
and_n #(2, 0, 0) AND_341 (fourFunc_wire_831, {fourFunc_wire_609_2, fourFunc_wire_610});
or_n #(2, 0, 0) OR_190 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_16_OR_intermediateXXXwire_690_AND_intermediateXXXwire_692, {NOT_intermediateXXXwire_690_AND_intermediateXXXwire_16, fourFunc_wire_831});
and_n #(2, 0, 0) AND_342 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_15, {fourFunc_wire_8_11, NOT_intermediateXXXwire_690_2});
and_n #(2, 0, 0) AND_343 (fourFunc_wire_832, {fourFunc_wire_609_3, fourFunc_wire_606});
or_n #(2, 0, 0) OR_191 (NOT_intermediateXXXwire_690_AND_intermediateXXXwire_15_OR_intermediateXXXwire_690_AND_intermediateXXXwire_688, {NOT_intermediateXXXwire_690_AND_intermediateXXXwire_15, fourFunc_wire_832});
and_n #(2, 0, 0) AND_344 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_757, {fourFunc_wire_552_1, NOT_intermediateXXXwire_697_0});
and_n #(2, 0, 0) AND_345 (fourFunc_wire_833, {fourFunc_wire_608_4, fourFunc_wire_745});
or_n #(2, 0, 0) OR_192 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_757_OR_intermediateXXXwire_697_AND_intermediateXXXwire_758, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_757, fourFunc_wire_833});
notg #(0, 0) NOT_119 (NOT_intermediateXXXwire_697, fourFunc_wire_608_5);
and_n #(2, 0, 0) AND_346 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_760, {fourFunc_wire_553_1, NOT_intermediateXXXwire_697_1});
and_n #(2, 0, 0) AND_347 (fourFunc_wire_834, {fourFunc_wire_608_6, fourFunc_wire_746});
or_n #(2, 0, 0) OR_193 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_760_OR_intermediateXXXwire_697_AND_intermediateXXXwire_761, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_760, fourFunc_wire_834});
and_n #(2, 0, 0) AND_348 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_763, {fourFunc_wire_554_1, NOT_intermediateXXXwire_697_2});
and_n #(2, 0, 0) AND_349 (fourFunc_wire_835, {fourFunc_wire_608_7, fourFunc_wire_747});
or_n #(2, 0, 0) OR_194 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_763_OR_intermediateXXXwire_697_AND_intermediateXXXwire_764, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_763, fourFunc_wire_835});
and_n #(2, 0, 0) AND_350 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_766, {fourFunc_wire_555_1, NOT_intermediateXXXwire_697_3});
and_n #(2, 0, 0) AND_351 (fourFunc_wire_836, {fourFunc_wire_608_8, fourFunc_wire_748});
or_n #(2, 0, 0) OR_195 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_766_OR_intermediateXXXwire_697_AND_intermediateXXXwire_767, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_766, fourFunc_wire_836});
and_n #(2, 0, 0) AND_352 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_769, {fourFunc_wire_556_1, NOT_intermediateXXXwire_697_4});
and_n #(2, 0, 0) AND_353 (fourFunc_wire_837, {fourFunc_wire_608_9, fourFunc_wire_749});
or_n #(2, 0, 0) OR_196 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_769_OR_intermediateXXXwire_697_AND_intermediateXXXwire_770, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_769, fourFunc_wire_837});
and_n #(2, 0, 0) AND_354 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_772, {fourFunc_wire_557_1, NOT_intermediateXXXwire_697_5});
and_n #(2, 0, 0) AND_355 (fourFunc_wire_838, {fourFunc_wire_608_10, fourFunc_wire_750});
or_n #(2, 0, 0) OR_197 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_772_OR_intermediateXXXwire_697_AND_intermediateXXXwire_773, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_772, fourFunc_wire_838});
and_n #(2, 0, 0) AND_356 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_775, {fourFunc_wire_558_1, NOT_intermediateXXXwire_697_6});
and_n #(2, 0, 0) AND_357 (fourFunc_wire_839, {fourFunc_wire_608_11, fourFunc_wire_751});
or_n #(2, 0, 0) OR_198 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_775_OR_intermediateXXXwire_697_AND_intermediateXXXwire_776, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_775, fourFunc_wire_839});
and_n #(2, 0, 0) AND_358 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_778, {fourFunc_wire_559_1, NOT_intermediateXXXwire_697_7});
and_n #(2, 0, 0) AND_359 (fourFunc_wire_840, {fourFunc_wire_608_12, fourFunc_wire_752});
or_n #(2, 0, 0) OR_199 (NOT_intermediateXXXwire_697_AND_intermediateXXXwire_778_OR_intermediateXXXwire_697_AND_intermediateXXXwire_779, {NOT_intermediateXXXwire_697_AND_intermediateXXXwire_778, fourFunc_wire_840});
and_n #(2, 0, 0) AND_360 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_914, {fourFunc_wire_53_18, NOT_intermediateXXXwire_922_0});
and_n #(2, 0, 0) AND_361 (fourFunc_wire_841, {fourFunc_wire_717_0, fourFunc_wire_809});
or_n #(2, 0, 0) OR_200 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_914_OR_intermediateXXXwire_922_AND_intermediateXXXwire_915, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_914, fourFunc_wire_841});
notg #(0, 0) NOT_120 (NOT_intermediateXXXwire_922, fourFunc_wire_717_1);
and_n #(2, 0, 0) AND_362 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_924, {fourFunc_wire_95_27, NOT_intermediateXXXwire_922_1});
and_n #(2, 0, 0) AND_363 (fourFunc_wire_842, {fourFunc_wire_717_2, fourFunc_wire_812});
or_n #(2, 0, 0) OR_201 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_924_OR_intermediateXXXwire_922_AND_intermediateXXXwire_925, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_924, fourFunc_wire_842});
and_n #(2, 0, 0) AND_364 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_932, {fourFunc_wire_90_14, NOT_intermediateXXXwire_922_2});
and_n #(2, 0, 0) AND_365 (fourFunc_wire_843, {fourFunc_wire_717_3, fourFunc_wire_814});
or_n #(2, 0, 0) OR_202 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_932_OR_intermediateXXXwire_922_AND_intermediateXXXwire_933, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_932, fourFunc_wire_843});
and_n #(2, 0, 0) AND_366 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_940, {fourFunc_wire_85_14, NOT_intermediateXXXwire_922_3});
and_n #(2, 0, 0) AND_367 (fourFunc_wire_844, {fourFunc_wire_717_4, fourFunc_wire_816});
or_n #(2, 0, 0) OR_203 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_940_OR_intermediateXXXwire_922_AND_intermediateXXXwire_941, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_940, fourFunc_wire_844});
and_n #(2, 0, 0) AND_368 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_948, {fourFunc_wire_80_14, NOT_intermediateXXXwire_922_4});
and_n #(2, 0, 0) AND_369 (fourFunc_wire_845, {fourFunc_wire_717_5, fourFunc_wire_818});
or_n #(2, 0, 0) OR_204 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_948_OR_intermediateXXXwire_922_AND_intermediateXXXwire_949, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_948, fourFunc_wire_845});
and_n #(2, 0, 0) AND_370 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_956, {fourFunc_wire_75_14, NOT_intermediateXXXwire_922_5});
and_n #(2, 0, 0) AND_371 (fourFunc_wire_846, {fourFunc_wire_717_6, fourFunc_wire_820});
or_n #(2, 0, 0) OR_205 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_956_OR_intermediateXXXwire_922_AND_intermediateXXXwire_957, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_956, fourFunc_wire_846});
and_n #(2, 0, 0) AND_372 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_964, {fourFunc_wire_70_14, NOT_intermediateXXXwire_922_6});
and_n #(2, 0, 0) AND_373 (fourFunc_wire_847, {fourFunc_wire_717_7, fourFunc_wire_822});
or_n #(2, 0, 0) OR_206 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_964_OR_intermediateXXXwire_922_AND_intermediateXXXwire_965, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_964, fourFunc_wire_847});
and_n #(2, 0, 0) AND_374 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_972, {fourFunc_wire_65_14, NOT_intermediateXXXwire_922_7});
and_n #(2, 0, 0) AND_375 (fourFunc_wire_848, {fourFunc_wire_717_8, fourFunc_wire_824});
or_n #(2, 0, 0) OR_207 (NOT_intermediateXXXwire_922_AND_intermediateXXXwire_972_OR_intermediateXXXwire_922_AND_intermediateXXXwire_973, {NOT_intermediateXXXwire_922_AND_intermediateXXXwire_972, fourFunc_wire_848});
and_n #(2, 0, 0) AND_376 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_781, {fourFunc_wire_54_5, NOT_intermediateXXXwire_795_0});
and_n #(2, 0, 0) AND_377 (fourFunc_wire_849, {fourFunc_wire_648_0, fourFunc_wire_753});
or_n #(2, 0, 0) OR_208 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_781_OR_intermediateXXXwire_795_AND_intermediateXXXwire_782, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_781, fourFunc_wire_849});
notg #(0, 0) NOT_121 (NOT_intermediateXXXwire_795, fourFunc_wire_648_1);
and_n #(2, 0, 0) AND_378 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_796, {fourFunc_wire_94_7, NOT_intermediateXXXwire_795_1});
and_n #(2, 0, 0) AND_379 (fourFunc_wire_850, {fourFunc_wire_648_2, fourFunc_wire_759});
or_n #(2, 0, 0) OR_209 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_796_OR_intermediateXXXwire_795_AND_intermediateXXXwire_797, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_796, fourFunc_wire_850});
and_n #(2, 0, 0) AND_380 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_809, {fourFunc_wire_89_7, NOT_intermediateXXXwire_795_2});
and_n #(2, 0, 0) AND_381 (fourFunc_wire_851, {fourFunc_wire_648_3, fourFunc_wire_765});
or_n #(2, 0, 0) OR_210 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_809_OR_intermediateXXXwire_795_AND_intermediateXXXwire_810, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_809, fourFunc_wire_851});
and_n #(2, 0, 0) AND_382 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_822, {fourFunc_wire_84_7, NOT_intermediateXXXwire_795_3});
and_n #(2, 0, 0) AND_383 (fourFunc_wire_852, {fourFunc_wire_648_4, fourFunc_wire_771});
or_n #(2, 0, 0) OR_211 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_822_OR_intermediateXXXwire_795_AND_intermediateXXXwire_823, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_822, fourFunc_wire_852});
and_n #(2, 0, 0) AND_384 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_835, {fourFunc_wire_79_7, NOT_intermediateXXXwire_795_4});
and_n #(2, 0, 0) AND_385 (fourFunc_wire_853, {fourFunc_wire_648_5, fourFunc_wire_777});
or_n #(2, 0, 0) OR_212 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_835_OR_intermediateXXXwire_795_AND_intermediateXXXwire_836, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_835, fourFunc_wire_853});
and_n #(2, 0, 0) AND_386 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_848, {fourFunc_wire_74_7, NOT_intermediateXXXwire_795_5});
and_n #(2, 0, 0) AND_387 (fourFunc_wire_854, {fourFunc_wire_648_6, fourFunc_wire_783});
or_n #(2, 0, 0) OR_213 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_848_OR_intermediateXXXwire_795_AND_intermediateXXXwire_849, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_848, fourFunc_wire_854});
and_n #(2, 0, 0) AND_388 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_861, {fourFunc_wire_69_7, NOT_intermediateXXXwire_795_6});
and_n #(2, 0, 0) AND_389 (fourFunc_wire_855, {fourFunc_wire_648_7, fourFunc_wire_789});
or_n #(2, 0, 0) OR_214 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_861_OR_intermediateXXXwire_795_AND_intermediateXXXwire_862, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_861, fourFunc_wire_855});
and_n #(2, 0, 0) AND_390 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_874, {fourFunc_wire_64_7, NOT_intermediateXXXwire_795_7});
and_n #(2, 0, 0) AND_391 (fourFunc_wire_856, {fourFunc_wire_648_8, fourFunc_wire_795});
or_n #(2, 0, 0) OR_215 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_874_OR_intermediateXXXwire_795_AND_intermediateXXXwire_875, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_874, fourFunc_wire_856});
and_n #(2, 0, 0) AND_392 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_887, {fourFunc_wire_59_5, NOT_intermediateXXXwire_795_8});
and_n #(2, 0, 0) AND_393 (fourFunc_wire_857, {fourFunc_wire_648_9, fourFunc_wire_801});
or_n #(2, 0, 0) OR_216 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_887_OR_intermediateXXXwire_795_AND_intermediateXXXwire_888, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_887, fourFunc_wire_857});
and_n #(2, 0, 0) AND_394 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_898, {fourFunc_wire_56_3, NOT_intermediateXXXwire_795_9});
and_n #(2, 0, 0) AND_395 (fourFunc_wire_858, {fourFunc_wire_648_10, fourFunc_wire_806});
or_n #(2, 0, 0) OR_217 (NOT_intermediateXXXwire_795_AND_intermediateXXXwire_898_OR_intermediateXXXwire_795_AND_intermediateXXXwire_899, {NOT_intermediateXXXwire_795_AND_intermediateXXXwire_898, fourFunc_wire_858});
dff DFF_1  (fourFunc_wire_551, NOT_intermediateXXXwire_676_AND_intermediateXXXwire_673_OR_intermediateXXXwire_676_AND_intermediateXXXwire_674, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_2  (fourFunc_wire_2, NOT_intermediateXXXwire_686_AND_intermediateXXXwire_14_OR_intermediateXXXwire_686_AND_intermediateXXXwire_682, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_3  (fourFunc_wire_10, NOT_intermediateXXXwire_690_AND_intermediateXXXwire_17_OR_intermediateXXXwire_690_AND_intermediateXXXwire_695, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_4  (fourFunc_wire_3, NOT_intermediateXXXwire_690_AND_intermediateXXXwire_16_OR_intermediateXXXwire_690_AND_intermediateXXXwire_692, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_5  (fourFunc_wire_8, NOT_intermediateXXXwire_690_AND_intermediateXXXwire_15_OR_intermediateXXXwire_690_AND_intermediateXXXwire_688, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_6  (fourFunc_wire_552, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_757_OR_intermediateXXXwire_697_AND_intermediateXXXwire_758, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_7  (fourFunc_wire_553, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_760_OR_intermediateXXXwire_697_AND_intermediateXXXwire_761, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_8  (fourFunc_wire_554, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_763_OR_intermediateXXXwire_697_AND_intermediateXXXwire_764, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_9  (fourFunc_wire_555, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_766_OR_intermediateXXXwire_697_AND_intermediateXXXwire_767, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_10  (fourFunc_wire_556, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_769_OR_intermediateXXXwire_697_AND_intermediateXXXwire_770, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_11  (fourFunc_wire_557, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_772_OR_intermediateXXXwire_697_AND_intermediateXXXwire_773, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_12  (fourFunc_wire_558, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_775_OR_intermediateXXXwire_697_AND_intermediateXXXwire_776, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_13  (fourFunc_wire_559, NOT_intermediateXXXwire_697_AND_intermediateXXXwire_778_OR_intermediateXXXwire_697_AND_intermediateXXXwire_779, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_14  (fourFunc_wire_53, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_914_OR_intermediateXXXwire_922_AND_intermediateXXXwire_915, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_15  (fourFunc_wire_95, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_924_OR_intermediateXXXwire_922_AND_intermediateXXXwire_925, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_16  (fourFunc_wire_90, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_932_OR_intermediateXXXwire_922_AND_intermediateXXXwire_933, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_17  (fourFunc_wire_85, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_940_OR_intermediateXXXwire_922_AND_intermediateXXXwire_941, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_18  (fourFunc_wire_80, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_948_OR_intermediateXXXwire_922_AND_intermediateXXXwire_949, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_19  (fourFunc_wire_75, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_956_OR_intermediateXXXwire_922_AND_intermediateXXXwire_957, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_20  (fourFunc_wire_70, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_964_OR_intermediateXXXwire_922_AND_intermediateXXXwire_965, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_21  (fourFunc_wire_65, NOT_intermediateXXXwire_922_AND_intermediateXXXwire_972_OR_intermediateXXXwire_922_AND_intermediateXXXwire_973, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_22  (fourFunc_wire_54, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_781_OR_intermediateXXXwire_795_AND_intermediateXXXwire_782, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_23  (fourFunc_wire_94, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_796_OR_intermediateXXXwire_795_AND_intermediateXXXwire_797, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_24  (fourFunc_wire_89, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_809_OR_intermediateXXXwire_795_AND_intermediateXXXwire_810, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_25  (fourFunc_wire_84, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_822_OR_intermediateXXXwire_795_AND_intermediateXXXwire_823, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_26  (fourFunc_wire_79, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_835_OR_intermediateXXXwire_795_AND_intermediateXXXwire_836, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_27  (fourFunc_wire_74, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_848_OR_intermediateXXXwire_795_AND_intermediateXXXwire_849, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_28  (fourFunc_wire_69, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_861_OR_intermediateXXXwire_795_AND_intermediateXXXwire_862, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_29  (fourFunc_wire_64, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_874_OR_intermediateXXXwire_795_AND_intermediateXXXwire_875, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_30  (fourFunc_wire_59, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_887_OR_intermediateXXXwire_795_AND_intermediateXXXwire_888, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_31  (fourFunc_wire_56, NOT_intermediateXXXwire_795_AND_intermediateXXXwire_898_OR_intermediateXXXwire_795_AND_intermediateXXXwire_899, fourFunc_wire_550, fourFunc_wire_549, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_32  (fourFunc_wire_592, fourFunc_wire_591, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_33  (fourFunc_wire_588, fourFunc_wire_593, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_34  (fourFunc_wire_589, fourFunc_wire_594, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_35  (fourFunc_wire_590, fourFunc_wire_595, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_36  (fourFunc_wire_586, fourFunc_wire_596, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_37  (fourFunc_wire_581, fourFunc_wire_597, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);
dff DFF_38  (fourFunc_wire_599, fourFunc_wire_598, fourFunc_wire_550, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0);

endmodule
